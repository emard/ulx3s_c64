);
end rom_kernal_pack;
