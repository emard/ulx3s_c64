);
end rom_chargen_pack;
