library IEEE;
use IEEE.std_logic_1164.all;

package rom_chargen_pack is
type t_rom_chargen is array(0 to 4095) of std_logic_vector(7 downto 0);
constant rom_chargen : t_rom_chargen :=
(
x"3C", x"66", x"6E", x"6E", x"60", x"66", x"3E", x"00",
x"3C", x"66", x"66", x"7E", x"66", x"66", x"66", x"00",
x"7C", x"66", x"66", x"7C", x"66", x"66", x"7E", x"00",
x"3C", x"66", x"66", x"60", x"60", x"66", x"3E", x"00",
x"7C", x"66", x"66", x"66", x"66", x"66", x"7C", x"00",
x"7E", x"66", x"60", x"78", x"60", x"66", x"7E", x"00",
x"7E", x"66", x"60", x"78", x"60", x"60", x"60", x"00",
x"3E", x"66", x"60", x"6E", x"66", x"66", x"3E", x"00",
x"66", x"66", x"66", x"7E", x"66", x"66", x"66", x"00",
x"7E", x"18", x"18", x"18", x"18", x"18", x"7E", x"00",
x"7E", x"66", x"06", x"06", x"66", x"66", x"7C", x"00",
x"66", x"66", x"6C", x"78", x"6C", x"66", x"66", x"00",
x"60", x"60", x"60", x"60", x"60", x"66", x"7E", x"00",
x"63", x"77", x"7F", x"7F", x"6B", x"63", x"63", x"00",
x"66", x"66", x"76", x"7E", x"6E", x"66", x"66", x"00",
x"3C", x"66", x"66", x"66", x"66", x"66", x"3E", x"00",
x"7C", x"66", x"66", x"7E", x"60", x"60", x"60", x"00",
x"3C", x"66", x"66", x"66", x"6A", x"6C", x"36", x"00",
x"7C", x"66", x"66", x"7C", x"66", x"66", x"66", x"00",
x"3E", x"60", x"70", x"3C", x"0E", x"0E", x"7C", x"00",
x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00",
x"66", x"66", x"66", x"66", x"66", x"6E", x"3C", x"00",
x"66", x"66", x"66", x"2C", x"3C", x"18", x"18", x"00",
x"63", x"63", x"6B", x"7F", x"7F", x"77", x"63", x"00",
x"66", x"66", x"3C", x"18", x"3C", x"66", x"66", x"00",
x"66", x"66", x"6E", x"3C", x"18", x"18", x"18", x"00",
x"7E", x"66", x"0C", x"18", x"30", x"76", x"7E", x"00",
x"3C", x"30", x"30", x"30", x"30", x"30", x"3C", x"00",
x"3C", x"66", x"60", x"78", x"30", x"30", x"7E", x"00",
x"3C", x"0C", x"0C", x"0C", x"0C", x"0C", x"3C", x"00",
x"08", x"1C", x"3E", x"1C", x"1C", x"1C", x"1C", x"00",
x"00", x"10", x"3F", x"7F", x"3F", x"10", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"38", x"38", x"38", x"38", x"38", x"00", x"38", x"00",
x"6C", x"6C", x"48", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"18", x"7E", x"60", x"7E", x"06", x"7E", x"18", x"00",
x"62", x"66", x"0C", x"18", x"30", x"66", x"46", x"00",
x"3C", x"66", x"66", x"3C", x"74", x"6E", x"3E", x"00",
x"18", x"18", x"10", x"00", x"00", x"00", x"00", x"00",
x"1C", x"30", x"30", x"30", x"30", x"30", x"1C", x"00",
x"38", x"0C", x"0C", x"0C", x"0C", x"0C", x"38", x"00",
x"08", x"2A", x"1C", x"7F", x"1C", x"2A", x"08", x"00",
x"00", x"18", x"18", x"7E", x"18", x"18", x"00", x"00",
x"00", x"00", x"00", x"00", x"18", x"18", x"08", x"00",
x"00", x"00", x"00", x"3C", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"00",
x"02", x"06", x"0C", x"18", x"30", x"60", x"40", x"00",
x"3C", x"66", x"6E", x"7E", x"76", x"66", x"3C", x"00",
x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00",
x"7C", x"66", x"06", x"1C", x"30", x"66", x"7E", x"00",
x"7C", x"66", x"06", x"0C", x"06", x"66", x"7E", x"00",
x"60", x"60", x"6C", x"7E", x"0C", x"0C", x"0C", x"00",
x"7E", x"66", x"60", x"7C", x"06", x"66", x"7C", x"00",
x"3E", x"66", x"60", x"7C", x"66", x"66", x"3E", x"00",
x"7E", x"66", x"06", x"1E", x"06", x"06", x"06", x"00",
x"3C", x"66", x"66", x"3C", x"66", x"66", x"7E", x"00",
x"3C", x"66", x"66", x"3E", x"06", x"66", x"7C", x"00",
x"00", x"18", x"18", x"00", x"18", x"18", x"00", x"00",
x"00", x"18", x"18", x"00", x"18", x"18", x"08", x"00",
x"00", x"0C", x"18", x"30", x"18", x"0C", x"00", x"00",
x"00", x"00", x"3C", x"00", x"3C", x"00", x"00", x"00",
x"00", x"30", x"18", x"0C", x"18", x"30", x"00", x"00",
x"7E", x"66", x"06", x"0C", x"18", x"00", x"18", x"00",
x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
x"08", x"1C", x"3E", x"7F", x"3E", x"1C", x"3E", x"00",
x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18",
x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00",
x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30",
x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C",
x"00", x"00", x"00", x"E0", x"F0", x"38", x"18", x"18",
x"18", x"18", x"1C", x"0F", x"07", x"00", x"00", x"00",
x"18", x"18", x"38", x"F0", x"E0", x"00", x"00", x"00",
x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"FF", x"FF",
x"C0", x"E0", x"70", x"38", x"1C", x"0E", x"07", x"03",
x"03", x"07", x"0E", x"1C", x"38", x"70", x"E0", x"C0",
x"FF", x"FF", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0",
x"FF", x"FF", x"03", x"03", x"03", x"03", x"03", x"03",
x"00", x"3C", x"7E", x"7E", x"7E", x"7E", x"3C", x"00",
x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00",
x"36", x"7F", x"7F", x"7F", x"3E", x"1C", x"08", x"00",
x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60",
x"00", x"00", x"00", x"07", x"0F", x"1C", x"18", x"18",
x"C3", x"E7", x"7E", x"3C", x"3C", x"7E", x"E7", x"C3",
x"00", x"3C", x"66", x"42", x"42", x"66", x"3C", x"00",
x"18", x"18", x"7E", x"7E", x"18", x"18", x"3C", x"00",
x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06",
x"08", x"1C", x"3E", x"7F", x"3E", x"1C", x"08", x"00",
x"18", x"18", x"18", x"FF", x"FF", x"18", x"18", x"18",
x"A0", x"50", x"A0", x"50", x"A0", x"50", x"A0", x"50",
x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18",
x"00", x"00", x"00", x"3E", x"76", x"36", x"36", x"00",
x"FF", x"7F", x"3F", x"1F", x"0F", x"07", x"03", x"01",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0",
x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0",
x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA", x"55",
x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03",
x"00", x"00", x"00", x"00", x"AA", x"55", x"AA", x"55",
x"FF", x"FE", x"FC", x"F8", x"F0", x"E0", x"C0", x"80",
x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03",
x"18", x"18", x"18", x"1F", x"1F", x"18", x"18", x"18",
x"00", x"00", x"00", x"00", x"0F", x"0F", x"0F", x"0F",
x"18", x"18", x"18", x"1F", x"1F", x"00", x"00", x"00",
x"00", x"00", x"00", x"F8", x"F8", x"18", x"18", x"18",
x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
x"00", x"00", x"00", x"1F", x"1F", x"18", x"18", x"18",
x"18", x"18", x"18", x"FF", x"FF", x"00", x"00", x"00",
x"00", x"00", x"00", x"FF", x"FF", x"18", x"18", x"18",
x"18", x"18", x"18", x"F8", x"F8", x"18", x"18", x"18",
x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0",
x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0",
x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07",
x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
x"03", x"03", x"03", x"03", x"03", x"03", x"FF", x"FF",
x"00", x"00", x"00", x"00", x"F0", x"F0", x"F0", x"F0",
x"0F", x"0F", x"0F", x"0F", x"00", x"00", x"00", x"00",
x"18", x"18", x"18", x"F8", x"F8", x"00", x"00", x"00",
x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"00", x"00",
x"F0", x"F0", x"F0", x"F0", x"0F", x"0F", x"0F", x"0F",
x"C3", x"99", x"91", x"91", x"9F", x"99", x"C1", x"FF",
x"C3", x"99", x"99", x"81", x"99", x"99", x"99", x"FF",
x"83", x"99", x"99", x"83", x"99", x"99", x"81", x"FF",
x"C3", x"99", x"99", x"9F", x"9F", x"99", x"C1", x"FF",
x"83", x"99", x"99", x"99", x"99", x"99", x"83", x"FF",
x"81", x"99", x"9F", x"87", x"9F", x"99", x"81", x"FF",
x"81", x"99", x"9F", x"87", x"9F", x"9F", x"9F", x"FF",
x"C1", x"99", x"9F", x"91", x"99", x"99", x"C1", x"FF",
x"99", x"99", x"99", x"81", x"99", x"99", x"99", x"FF",
x"81", x"E7", x"E7", x"E7", x"E7", x"E7", x"81", x"FF",
x"81", x"99", x"F9", x"F9", x"99", x"99", x"83", x"FF",
x"99", x"99", x"93", x"87", x"93", x"99", x"99", x"FF",
x"9F", x"9F", x"9F", x"9F", x"9F", x"99", x"81", x"FF",
x"9C", x"88", x"80", x"80", x"94", x"9C", x"9C", x"FF",
x"99", x"99", x"89", x"81", x"91", x"99", x"99", x"FF",
x"C3", x"99", x"99", x"99", x"99", x"99", x"C1", x"FF",
x"83", x"99", x"99", x"81", x"9F", x"9F", x"9F", x"FF",
x"C3", x"99", x"99", x"99", x"95", x"93", x"C9", x"FF",
x"83", x"99", x"99", x"83", x"99", x"99", x"99", x"FF",
x"C1", x"9F", x"8F", x"C3", x"F1", x"F1", x"83", x"FF",
x"81", x"E7", x"E7", x"E7", x"E7", x"E7", x"E7", x"FF",
x"99", x"99", x"99", x"99", x"99", x"91", x"C3", x"FF",
x"99", x"99", x"99", x"D3", x"C3", x"E7", x"E7", x"FF",
x"9C", x"9C", x"94", x"80", x"80", x"88", x"9C", x"FF",
x"99", x"99", x"C3", x"E7", x"C3", x"99", x"99", x"FF",
x"99", x"99", x"91", x"C3", x"E7", x"E7", x"E7", x"FF",
x"81", x"99", x"F3", x"E7", x"CF", x"89", x"81", x"FF",
x"C3", x"CF", x"CF", x"CF", x"CF", x"CF", x"C3", x"FF",
x"C3", x"99", x"9F", x"87", x"CF", x"CF", x"81", x"FF",
x"C3", x"F3", x"F3", x"F3", x"F3", x"F3", x"C3", x"FF",
x"F7", x"E3", x"C1", x"E3", x"E3", x"E3", x"E3", x"FF",
x"FF", x"EF", x"C0", x"80", x"C0", x"EF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"C7", x"C7", x"C7", x"C7", x"C7", x"FF", x"C7", x"FF",
x"93", x"93", x"B7", x"FF", x"FF", x"FF", x"FF", x"FF",
x"C9", x"C9", x"80", x"C9", x"80", x"C9", x"C9", x"FF",
x"E7", x"81", x"9F", x"81", x"F9", x"81", x"E7", x"FF",
x"9D", x"99", x"F3", x"E7", x"CF", x"99", x"B9", x"FF",
x"C3", x"99", x"99", x"C3", x"8B", x"91", x"C1", x"FF",
x"E7", x"E7", x"EF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"E3", x"CF", x"CF", x"CF", x"CF", x"CF", x"E3", x"FF",
x"C7", x"F3", x"F3", x"F3", x"F3", x"F3", x"C7", x"FF",
x"F7", x"D5", x"E3", x"80", x"E3", x"D5", x"F7", x"FF",
x"FF", x"E7", x"E7", x"81", x"E7", x"E7", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"E7", x"E7", x"F7", x"FF",
x"FF", x"FF", x"FF", x"C3", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"E7", x"E7", x"FF",
x"FD", x"F9", x"F3", x"E7", x"CF", x"9F", x"BF", x"FF",
x"C3", x"99", x"91", x"81", x"89", x"99", x"C3", x"FF",
x"E7", x"C7", x"E7", x"E7", x"E7", x"E7", x"81", x"FF",
x"83", x"99", x"F9", x"E3", x"CF", x"99", x"81", x"FF",
x"83", x"99", x"F9", x"F3", x"F9", x"99", x"81", x"FF",
x"9F", x"9F", x"93", x"81", x"F3", x"F3", x"F3", x"FF",
x"81", x"99", x"9F", x"83", x"F9", x"99", x"83", x"FF",
x"C1", x"99", x"9F", x"83", x"99", x"99", x"C1", x"FF",
x"81", x"99", x"F9", x"E1", x"F9", x"F9", x"F9", x"FF",
x"C3", x"99", x"99", x"C3", x"99", x"99", x"81", x"FF",
x"C3", x"99", x"99", x"C1", x"F9", x"99", x"83", x"FF",
x"FF", x"E7", x"E7", x"FF", x"E7", x"E7", x"FF", x"FF",
x"FF", x"E7", x"E7", x"FF", x"E7", x"E7", x"F7", x"FF",
x"FF", x"F3", x"E7", x"CF", x"E7", x"F3", x"FF", x"FF",
x"FF", x"FF", x"C3", x"FF", x"C3", x"FF", x"FF", x"FF",
x"FF", x"CF", x"E7", x"F3", x"E7", x"CF", x"FF", x"FF",
x"81", x"99", x"F9", x"F3", x"E7", x"FF", x"E7", x"FF",
x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
x"F7", x"E3", x"C1", x"80", x"C1", x"E3", x"C1", x"FF",
x"E7", x"E7", x"E7", x"E7", x"E7", x"E7", x"E7", x"E7",
x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
x"CF", x"CF", x"CF", x"CF", x"CF", x"CF", x"CF", x"CF",
x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3",
x"FF", x"FF", x"FF", x"1F", x"0F", x"C7", x"E7", x"E7",
x"E7", x"E7", x"E3", x"F0", x"F8", x"FF", x"FF", x"FF",
x"E7", x"E7", x"C7", x"0F", x"1F", x"FF", x"FF", x"FF",
x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"00", x"00",
x"3F", x"1F", x"8F", x"C7", x"E3", x"F1", x"F8", x"FC",
x"FC", x"F8", x"F1", x"E3", x"C7", x"8F", x"1F", x"3F",
x"00", x"00", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F",
x"00", x"00", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
x"FF", x"C3", x"81", x"81", x"81", x"81", x"C3", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
x"C9", x"80", x"80", x"80", x"C1", x"E3", x"F7", x"FF",
x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F",
x"FF", x"FF", x"FF", x"F8", x"F0", x"E3", x"E7", x"E7",
x"3C", x"18", x"81", x"C3", x"C3", x"81", x"18", x"3C",
x"FF", x"C3", x"99", x"BD", x"BD", x"99", x"C3", x"FF",
x"E7", x"E7", x"81", x"81", x"E7", x"E7", x"C3", x"FF",
x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9",
x"F7", x"E3", x"C1", x"80", x"C1", x"E3", x"F7", x"FF",
x"E7", x"E7", x"E7", x"00", x"00", x"E7", x"E7", x"E7",
x"5F", x"AF", x"5F", x"AF", x"5F", x"AF", x"5F", x"AF",
x"E7", x"E7", x"E7", x"E7", x"E7", x"E7", x"E7", x"E7",
x"FF", x"FF", x"FF", x"C1", x"89", x"C9", x"C9", x"FF",
x"00", x"80", x"C0", x"E0", x"F0", x"F8", x"FC", x"FE",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F",
x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F",
x"55", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA",
x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
x"FF", x"FF", x"FF", x"FF", x"55", x"AA", x"55", x"AA",
x"00", x"01", x"03", x"07", x"0F", x"1F", x"3F", x"7F",
x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
x"E7", x"E7", x"E7", x"E0", x"E0", x"E7", x"E7", x"E7",
x"FF", x"FF", x"FF", x"FF", x"F0", x"F0", x"F0", x"F0",
x"E7", x"E7", x"E7", x"E0", x"E0", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"07", x"07", x"E7", x"E7", x"E7",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
x"FF", x"FF", x"FF", x"E0", x"E0", x"E7", x"E7", x"E7",
x"E7", x"E7", x"E7", x"00", x"00", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"00", x"00", x"E7", x"E7", x"E7",
x"E7", x"E7", x"E7", x"07", x"07", x"E7", x"E7", x"E7",
x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F",
x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F",
x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8",
x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"00", x"00",
x"FF", x"FF", x"FF", x"FF", x"0F", x"0F", x"0F", x"0F",
x"F0", x"F0", x"F0", x"F0", x"FF", x"FF", x"FF", x"FF",
x"E7", x"E7", x"E7", x"07", x"07", x"FF", x"FF", x"FF",
x"0F", x"0F", x"0F", x"0F", x"FF", x"FF", x"FF", x"FF",
x"0F", x"0F", x"0F", x"0F", x"F0", x"F0", x"F0", x"F0",
x"3C", x"66", x"6E", x"6E", x"60", x"66", x"3E", x"00",
x"00", x"00", x"3C", x"06", x"3E", x"66", x"7E", x"00",
x"00", x"60", x"60", x"7C", x"66", x"66", x"7E", x"00",
x"00", x"00", x"3E", x"60", x"60", x"60", x"7E", x"00",
x"00", x"06", x"06", x"3E", x"66", x"66", x"7E", x"00",
x"00", x"00", x"3C", x"66", x"7E", x"60", x"7E", x"00",
x"00", x"0E", x"18", x"3C", x"18", x"18", x"18", x"00",
x"00", x"00", x"3E", x"66", x"66", x"7E", x"06", x"3C",
x"00", x"60", x"60", x"7C", x"66", x"66", x"66", x"00",
x"00", x"18", x"00", x"18", x"18", x"18", x"18", x"00",
x"00", x"0C", x"00", x"0C", x"0C", x"0C", x"6C", x"78",
x"00", x"60", x"66", x"6C", x"78", x"6C", x"66", x"00",
x"00", x"18", x"18", x"18", x"18", x"18", x"3C", x"00",
x"00", x"00", x"7E", x"6B", x"6B", x"63", x"63", x"00",
x"00", x"00", x"7C", x"66", x"66", x"66", x"66", x"00",
x"00", x"00", x"3C", x"66", x"66", x"66", x"3E", x"00",
x"00", x"00", x"7C", x"66", x"66", x"7E", x"60", x"60",
x"00", x"00", x"3E", x"66", x"66", x"7E", x"06", x"06",
x"00", x"00", x"7E", x"66", x"60", x"60", x"60", x"00",
x"00", x"00", x"3E", x"60", x"7E", x"06", x"7E", x"00",
x"00", x"18", x"7E", x"18", x"18", x"18", x"1C", x"00",
x"00", x"00", x"66", x"66", x"66", x"66", x"3E", x"00",
x"00", x"00", x"66", x"66", x"66", x"34", x"18", x"00",
x"00", x"00", x"63", x"63", x"6B", x"6B", x"3F", x"00",
x"00", x"00", x"66", x"3C", x"18", x"3C", x"66", x"00",
x"00", x"00", x"66", x"66", x"66", x"3C", x"18", x"30",
x"00", x"00", x"7E", x"0C", x"18", x"30", x"7E", x"00",
x"3C", x"30", x"30", x"30", x"30", x"30", x"3C", x"00",
x"3C", x"66", x"60", x"78", x"30", x"30", x"7E", x"00",
x"3C", x"0C", x"0C", x"0C", x"0C", x"0C", x"3C", x"00",
x"08", x"1C", x"3E", x"1C", x"1C", x"1C", x"1C", x"00",
x"00", x"10", x"3F", x"7F", x"3F", x"10", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"38", x"38", x"38", x"38", x"38", x"00", x"38", x"00",
x"6C", x"6C", x"48", x"00", x"00", x"00", x"00", x"00",
x"36", x"36", x"7F", x"36", x"7F", x"36", x"36", x"00",
x"18", x"7E", x"60", x"7E", x"06", x"7E", x"18", x"00",
x"62", x"66", x"0C", x"18", x"30", x"66", x"46", x"00",
x"3C", x"66", x"66", x"3C", x"74", x"6E", x"3E", x"00",
x"18", x"18", x"10", x"00", x"00", x"00", x"00", x"00",
x"1C", x"30", x"30", x"30", x"30", x"30", x"1C", x"00",
x"38", x"0C", x"0C", x"0C", x"0C", x"0C", x"38", x"00",
x"08", x"2A", x"1C", x"7F", x"1C", x"2A", x"08", x"00",
x"00", x"18", x"18", x"7E", x"18", x"18", x"00", x"00",
x"00", x"00", x"00", x"00", x"18", x"18", x"08", x"00",
x"00", x"00", x"00", x"3C", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"00",
x"02", x"06", x"0C", x"18", x"30", x"60", x"40", x"00",
x"3C", x"66", x"6E", x"7E", x"76", x"66", x"3C", x"00",
x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00",
x"7C", x"66", x"06", x"1C", x"30", x"66", x"7E", x"00",
x"7C", x"66", x"06", x"0C", x"06", x"66", x"7E", x"00",
x"60", x"60", x"6C", x"7E", x"0C", x"0C", x"0C", x"00",
x"7E", x"66", x"60", x"7C", x"06", x"66", x"7C", x"00",
x"3E", x"66", x"60", x"7C", x"66", x"66", x"3E", x"00",
x"7E", x"66", x"06", x"1E", x"06", x"06", x"06", x"00",
x"3C", x"66", x"66", x"3C", x"66", x"66", x"7E", x"00",
x"3C", x"66", x"66", x"3E", x"06", x"66", x"7C", x"00",
x"00", x"18", x"18", x"00", x"18", x"18", x"00", x"00",
x"00", x"18", x"18", x"00", x"18", x"18", x"08", x"00",
x"00", x"0C", x"18", x"30", x"18", x"0C", x"00", x"00",
x"00", x"00", x"3C", x"00", x"3C", x"00", x"00", x"00",
x"00", x"30", x"18", x"0C", x"18", x"30", x"00", x"00",
x"7E", x"66", x"06", x"0C", x"18", x"00", x"18", x"00",
x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
x"3C", x"66", x"66", x"7E", x"66", x"66", x"66", x"00",
x"7C", x"66", x"66", x"7C", x"66", x"66", x"7E", x"00",
x"3C", x"66", x"66", x"60", x"60", x"66", x"3E", x"00",
x"7C", x"66", x"66", x"66", x"66", x"66", x"7C", x"00",
x"7E", x"66", x"60", x"78", x"60", x"66", x"7E", x"00",
x"7E", x"66", x"60", x"78", x"60", x"60", x"60", x"00",
x"3E", x"66", x"60", x"6E", x"66", x"66", x"3E", x"00",
x"66", x"66", x"66", x"7E", x"66", x"66", x"66", x"00",
x"7E", x"18", x"18", x"18", x"18", x"18", x"7E", x"00",
x"7E", x"66", x"06", x"06", x"66", x"66", x"7C", x"00",
x"66", x"66", x"6C", x"78", x"6C", x"66", x"66", x"00",
x"60", x"60", x"60", x"60", x"60", x"66", x"7E", x"00",
x"63", x"77", x"7F", x"7F", x"6B", x"63", x"63", x"00",
x"66", x"66", x"76", x"7E", x"6E", x"66", x"66", x"00",
x"3C", x"66", x"66", x"66", x"66", x"66", x"3E", x"00",
x"7C", x"66", x"66", x"7E", x"60", x"60", x"60", x"00",
x"3C", x"66", x"66", x"66", x"6A", x"6C", x"36", x"00",
x"7C", x"66", x"66", x"7C", x"66", x"66", x"66", x"00",
x"3E", x"60", x"70", x"3C", x"0E", x"0E", x"7C", x"00",
x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00",
x"66", x"66", x"66", x"66", x"66", x"6E", x"3C", x"00",
x"66", x"66", x"66", x"2C", x"3C", x"18", x"18", x"00",
x"63", x"63", x"6B", x"7F", x"7F", x"77", x"63", x"00",
x"66", x"66", x"3C", x"18", x"3C", x"66", x"66", x"00",
x"66", x"66", x"6E", x"3C", x"18", x"18", x"18", x"00",
x"7E", x"66", x"0C", x"18", x"30", x"76", x"7E", x"00",
x"18", x"18", x"18", x"FF", x"FF", x"18", x"18", x"18",
x"C0", x"C0", x"30", x"30", x"C0", x"C0", x"30", x"30",
x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18",
x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA", x"55",
x"33", x"99", x"CC", x"66", x"33", x"99", x"CC", x"66",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0",
x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0",
x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA", x"55",
x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03",
x"00", x"00", x"00", x"00", x"AA", x"55", x"AA", x"55",
x"CC", x"99", x"33", x"66", x"CC", x"99", x"33", x"66",
x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03",
x"18", x"18", x"18", x"1F", x"1F", x"18", x"18", x"18",
x"00", x"00", x"00", x"00", x"0F", x"0F", x"0F", x"0F",
x"18", x"18", x"18", x"1F", x"1F", x"00", x"00", x"00",
x"00", x"00", x"00", x"F8", x"F8", x"18", x"18", x"18",
x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
x"00", x"00", x"00", x"1F", x"1F", x"18", x"18", x"18",
x"18", x"18", x"18", x"FF", x"FF", x"00", x"00", x"00",
x"00", x"00", x"00", x"FF", x"FF", x"18", x"18", x"18",
x"18", x"18", x"18", x"F8", x"F8", x"18", x"18", x"18",
x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0",
x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0",
x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07",
x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
x"00", x"01", x"03", x"46", x"6C", x"38", x"10", x"00",
x"00", x"00", x"00", x"00", x"F0", x"F0", x"F0", x"F0",
x"0F", x"0F", x"0F", x"0F", x"00", x"00", x"00", x"00",
x"18", x"18", x"18", x"F8", x"F8", x"00", x"00", x"00",
x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"00", x"00",
x"F0", x"F0", x"F0", x"F0", x"0F", x"0F", x"0F", x"0F",
x"C3", x"99", x"91", x"91", x"9F", x"99", x"C1", x"FF",
x"FF", x"FF", x"C3", x"F9", x"C1", x"99", x"81", x"FF",
x"FF", x"9F", x"9F", x"83", x"99", x"99", x"81", x"FF",
x"FF", x"FF", x"C1", x"9F", x"9F", x"9F", x"81", x"FF",
x"FF", x"F9", x"F9", x"C1", x"99", x"99", x"81", x"FF",
x"FF", x"FF", x"C3", x"99", x"81", x"9F", x"81", x"FF",
x"FF", x"F1", x"E7", x"C3", x"E7", x"E7", x"E7", x"FF",
x"FF", x"FF", x"C1", x"99", x"99", x"81", x"F9", x"C3",
x"FF", x"9F", x"9F", x"83", x"99", x"99", x"99", x"FF",
x"FF", x"E7", x"FF", x"E7", x"E7", x"E7", x"E7", x"FF",
x"FF", x"F3", x"FF", x"F3", x"F3", x"F3", x"93", x"87",
x"FF", x"9F", x"99", x"93", x"87", x"93", x"99", x"FF",
x"FF", x"E7", x"E7", x"E7", x"E7", x"E7", x"C3", x"FF",
x"FF", x"FF", x"81", x"94", x"94", x"9C", x"9C", x"FF",
x"FF", x"FF", x"83", x"99", x"99", x"99", x"99", x"FF",
x"FF", x"FF", x"C3", x"99", x"99", x"99", x"C1", x"FF",
x"FF", x"FF", x"83", x"99", x"99", x"81", x"9F", x"9F",
x"FF", x"FF", x"C1", x"99", x"99", x"81", x"F9", x"F9",
x"FF", x"FF", x"81", x"99", x"9F", x"9F", x"9F", x"FF",
x"FF", x"FF", x"C1", x"9F", x"81", x"F9", x"81", x"FF",
x"FF", x"E7", x"81", x"E7", x"E7", x"E7", x"E3", x"FF",
x"FF", x"FF", x"99", x"99", x"99", x"99", x"C1", x"FF",
x"FF", x"FF", x"99", x"99", x"99", x"CB", x"E7", x"FF",
x"FF", x"FF", x"9C", x"9C", x"94", x"94", x"C0", x"FF",
x"FF", x"FF", x"99", x"C3", x"E7", x"C3", x"99", x"FF",
x"FF", x"FF", x"99", x"99", x"99", x"C3", x"E7", x"CF",
x"FF", x"FF", x"81", x"F3", x"E7", x"CF", x"81", x"FF",
x"C3", x"CF", x"CF", x"CF", x"CF", x"CF", x"C3", x"FF",
x"C3", x"99", x"9F", x"87", x"CF", x"CF", x"81", x"FF",
x"C3", x"F3", x"F3", x"F3", x"F3", x"F3", x"C3", x"FF",
x"F7", x"E3", x"C1", x"E3", x"E3", x"E3", x"E3", x"FF",
x"FF", x"EF", x"C0", x"80", x"C0", x"EF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"C7", x"C7", x"C7", x"C7", x"C7", x"FF", x"C7", x"FF",
x"93", x"93", x"B7", x"FF", x"FF", x"FF", x"FF", x"FF",
x"C9", x"C9", x"80", x"C9", x"80", x"C9", x"C9", x"FF",
x"E7", x"81", x"9F", x"81", x"F9", x"81", x"E7", x"FF",
x"9D", x"99", x"F3", x"E7", x"CF", x"99", x"B9", x"FF",
x"C3", x"99", x"99", x"C3", x"8B", x"91", x"C1", x"FF",
x"E7", x"E7", x"EF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"E3", x"CF", x"CF", x"CF", x"CF", x"CF", x"E3", x"FF",
x"C7", x"F3", x"F3", x"F3", x"F3", x"F3", x"C7", x"FF",
x"F7", x"D5", x"E3", x"80", x"E3", x"D5", x"F7", x"FF",
x"FF", x"E7", x"E7", x"81", x"E7", x"E7", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"E7", x"E7", x"F7", x"FF",
x"FF", x"FF", x"FF", x"C3", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"E7", x"E7", x"FF",
x"FD", x"F9", x"F3", x"E7", x"CF", x"9F", x"BF", x"FF",
x"C3", x"99", x"91", x"81", x"89", x"99", x"C3", x"FF",
x"E7", x"C7", x"E7", x"E7", x"E7", x"E7", x"81", x"FF",
x"83", x"99", x"F9", x"E3", x"CF", x"99", x"81", x"FF",
x"83", x"99", x"F9", x"F3", x"F9", x"99", x"81", x"FF",
x"9F", x"9F", x"93", x"81", x"F3", x"F3", x"F3", x"FF",
x"81", x"99", x"9F", x"83", x"F9", x"99", x"83", x"FF",
x"C1", x"99", x"9F", x"83", x"99", x"99", x"C1", x"FF",
x"81", x"99", x"F9", x"E1", x"F9", x"F9", x"F9", x"FF",
x"C3", x"99", x"99", x"C3", x"99", x"99", x"81", x"FF",
x"C3", x"99", x"99", x"C1", x"F9", x"99", x"83", x"FF",
x"FF", x"E7", x"E7", x"FF", x"E7", x"E7", x"FF", x"FF",
x"FF", x"E7", x"E7", x"FF", x"E7", x"E7", x"F7", x"FF",
x"FF", x"F3", x"E7", x"CF", x"E7", x"F3", x"FF", x"FF",
x"FF", x"FF", x"C3", x"FF", x"C3", x"FF", x"FF", x"FF",
x"FF", x"CF", x"E7", x"F3", x"E7", x"CF", x"FF", x"FF",
x"81", x"99", x"F9", x"F3", x"E7", x"FF", x"E7", x"FF",
x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
x"C3", x"99", x"99", x"81", x"99", x"99", x"99", x"FF",
x"83", x"99", x"99", x"83", x"99", x"99", x"81", x"FF",
x"C3", x"99", x"99", x"9F", x"9F", x"99", x"C1", x"FF",
x"83", x"99", x"99", x"99", x"99", x"99", x"83", x"FF",
x"81", x"99", x"9F", x"87", x"9F", x"99", x"81", x"FF",
x"81", x"99", x"9F", x"87", x"9F", x"9F", x"9F", x"FF",
x"C1", x"99", x"9F", x"91", x"99", x"99", x"C1", x"FF",
x"99", x"99", x"99", x"81", x"99", x"99", x"99", x"FF",
x"81", x"E7", x"E7", x"E7", x"E7", x"E7", x"81", x"FF",
x"81", x"99", x"F9", x"F9", x"99", x"99", x"83", x"FF",
x"99", x"99", x"93", x"87", x"93", x"99", x"99", x"FF",
x"9F", x"9F", x"9F", x"9F", x"9F", x"99", x"81", x"FF",
x"9C", x"88", x"80", x"80", x"94", x"9C", x"9C", x"FF",
x"99", x"99", x"89", x"81", x"91", x"99", x"99", x"FF",
x"C3", x"99", x"99", x"99", x"99", x"99", x"C1", x"FF",
x"83", x"99", x"99", x"81", x"9F", x"9F", x"9F", x"FF",
x"C3", x"99", x"99", x"99", x"95", x"93", x"C9", x"FF",
x"83", x"99", x"99", x"83", x"99", x"99", x"99", x"FF",
x"C1", x"9F", x"8F", x"C3", x"F1", x"F1", x"83", x"FF",
x"81", x"E7", x"E7", x"E7", x"E7", x"E7", x"E7", x"FF",
x"99", x"99", x"99", x"99", x"99", x"91", x"C3", x"FF",
x"99", x"99", x"99", x"D3", x"C3", x"E7", x"E7", x"FF",
x"9C", x"9C", x"94", x"80", x"80", x"88", x"9C", x"FF",
x"99", x"99", x"C3", x"E7", x"C3", x"99", x"99", x"FF",
x"99", x"99", x"91", x"C3", x"E7", x"E7", x"E7", x"FF",
x"81", x"99", x"F3", x"E7", x"CF", x"89", x"81", x"FF",
x"E7", x"E7", x"E7", x"00", x"00", x"E7", x"E7", x"E7",
x"3F", x"3F", x"CF", x"CF", x"3F", x"3F", x"CF", x"CF",
x"E7", x"E7", x"E7", x"E7", x"E7", x"E7", x"E7", x"E7",
x"55", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA",
x"CC", x"66", x"33", x"99", x"CC", x"66", x"33", x"99",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F",
x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F",
x"55", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA",
x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
x"FF", x"FF", x"FF", x"FF", x"55", x"AA", x"55", x"AA",
x"33", x"66", x"CC", x"99", x"33", x"66", x"CC", x"99",
x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
x"E7", x"E7", x"E7", x"E0", x"E0", x"E7", x"E7", x"E7",
x"FF", x"FF", x"FF", x"FF", x"F0", x"F0", x"F0", x"F0",
x"E7", x"E7", x"E7", x"E0", x"E0", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"07", x"07", x"E7", x"E7", x"E7",
x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
x"FF", x"FF", x"FF", x"E0", x"E0", x"E7", x"E7", x"E7",
x"E7", x"E7", x"E7", x"00", x"00", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"00", x"00", x"E7", x"E7", x"E7",
x"E7", x"E7", x"E7", x"07", x"07", x"E7", x"E7", x"E7",
x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F",
x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F",
x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8",
x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
x"FF", x"FE", x"FC", x"B9", x"93", x"C7", x"EF", x"FF",
x"FF", x"FF", x"FF", x"FF", x"0F", x"0F", x"0F", x"0F",
x"F0", x"F0", x"F0", x"F0", x"FF", x"FF", x"FF", x"FF",
x"E7", x"E7", x"E7", x"07", x"07", x"FF", x"FF", x"FF",
x"0F", x"0F", x"0F", x"0F", x"FF", x"FF", x"FF", x"FF",
x"0F", x"0F", x"0F", x"0F", x"F0", x"F0", x"F0", x"F0"
);
end rom_chargen_pack;
