library IEEE;
use IEEE.std_logic_1164.all;

package rom_kernal_pack is
type t_rom_kernal is array(0 to 16383) of std_logic_vector(7 downto 0);
constant rom_kernal : t_rom_kernal :=
(
x"94", x"E3", x"B7", x"E3", x"4F", x"52", x"47", x"42",
x"41", x"53", x"49", x"43", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"A0", x"00", x"20",
x"88", x"E1", x"E6", x"7A", x"D0", x"02", x"E6", x"7B",
x"60", x"8B", x"E3", x"83", x"A4", x"7C", x"A5", x"1A",
x"A7", x"E4", x"A7", x"86", x"AE", x"8F", x"BA", x"A5",
x"BB", x"20", x"76", x"A1", x"B0", x"01", x"60", x"C9",
x"30", x"90", x"0A", x"C9", x"3A", x"60", x"C9", x"41",
x"90", x"03", x"C9", x"7B", x"60", x"38", x"60", x"20",
x"45", x"BC", x"20", x"4D", x"A1", x"20", x"4D", x"A1",
x"C9", x"4C", x"F0", x"03", x"4C", x"CF", x"A6", x"20",
x"E1", x"B3", x"4C", x"B3", x"BA", x"A9", x"00", x"85",
x"26", x"85", x"27", x"85", x"28", x"85", x"29", x"85",
x"2A", x"60", x"18", x"65", x"26", x"85", x"26", x"90",
x"02", x"E6", x"27", x"60", x"A5", x"62", x"85", x"8F",
x"45", x"63", x"85", x"8E", x"45", x"64", x"85", x"8D",
x"45", x"65", x"85", x"8C", x"45", x"61", x"85", x"8B",
x"4C", x"BE", x"E0", x"20", x"1B", x"A7", x"B0", x"11",
x"A9", x"0D", x"20", x"2E", x"BA", x"B0", x"0A", x"A5",
x"15", x"F0", x"03", x"4C", x"CC", x"A6", x"A5", x"14",
x"18", x"60", x"20", x"60", x"E0", x"20", x"7F", x"AF",
x"C9", x"3A", x"D0", x"03", x"4C", x"93", x"A4", x"C9",
x"00", x"D0", x"03", x"4C", x"E9", x"A4", x"4C", x"CF",
x"A6", x"A5", x"B0", x"05", x"B1", x"F0", x"0F", x"A2",
x"06", x"20", x"59", x"B9", x"A5", x"B1", x"20", x"0D",
x"FB", x"A5", x"B0", x"20", x"0D", x"FB", x"4C", x"34",
x"AC", x"85", x"50", x"38", x"A5", x"33", x"E5", x"50",
x"85", x"33", x"B0", x"02", x"C6", x"34", x"A5", x"32",
x"C5", x"34", x"F0", x"01", x"60", x"A5", x"31", x"C5",
x"33", x"60", x"4D", x"04", x"DC", x"85", x"8E", x"8A",
x"4D", x"12", x"D0", x"85", x"8C", x"98", x"4D", x"05",
x"DC", x"85", x"8F", x"A5", x"A2", x"4D", x"1B", x"D4",
x"85", x"8D", x"4C", x"BE", x"E0", x"84", x"2A", x"38",
x"A5", x"24", x"E5", x"2A", x"85", x"24", x"B0", x"02",
x"C6", x"25", x"38", x"A5", x"26", x"E5", x"2A", x"85",
x"26", x"B0", x"02", x"C6", x"27", x"E6", x"29", x"60",
x"3E", x"3D", x"3C", x"2F", x"2D", x"2A", x"5E", x"2B",
x"51", x"23", x"28", x"4B", x"58", x"59", x"57", x"48",
x"56", x"42", x"4D", x"24", x"47", x"43", x"0D", x"27",
x"5A", x"2E", x"4A", x"3F", x"20", x"1E", x"BC", x"20",
x"2E", x"BA", x"B0", x"0B", x"20", x"7F", x"AF", x"C9",
x"2C", x"F0", x"07", x"C9", x"29", x"F0", x"06", x"4C",
x"CF", x"A6", x"A0", x"00", x"60", x"A0", x"FF", x"60",
x"20", x"D2", x"F7", x"A2", x"1D", x"20", x"53", x"B9",
x"A5", x"3A", x"C9", x"FF", x"F0", x"0C", x"A2", x"04",
x"20", x"59", x"B9", x"A5", x"3A", x"A6", x"39", x"20",
x"51", x"B4", x"4C", x"32", x"AC", x"A5", x"6D", x"85",
x"65", x"A5", x"6C", x"85", x"64", x"A5", x"6B", x"85",
x"63", x"A5", x"6A", x"85", x"62", x"A5", x"6E", x"85",
x"66", x"A5", x"69", x"85", x"61", x"A2", x"00", x"86",
x"70", x"60", x"A5", x"61", x"F0", x"22", x"A5", x"70",
x"10", x"1A", x"E6", x"65", x"D0", x"16", x"E6", x"64",
x"D0", x"12", x"E6", x"63", x"D0", x"0E", x"E6", x"62",
x"D0", x"0A", x"A9", x"80", x"85", x"62", x"E6", x"61",
x"D0", x"02", x"C6", x"61", x"A9", x"00", x"85", x"70",
x"60", x"A0", x"00", x"20", x"95", x"E1", x"85", x"0B",
x"C8", x"20", x"95", x"E1", x"85", x"0F", x"A5", x"0B",
x"38", x"E5", x"3D", x"85", x"0B", x"A5", x"0F", x"E5",
x"3E", x"85", x"0F", x"A5", x"0F", x"E9", x"00", x"C9",
x"00", x"F0", x"03", x"4C", x"B0", x"A6", x"A6", x"0B",
x"20", x"C4", x"BF", x"4C", x"DE", x"A7", x"A9", x"01",
x"85", x"2B", x"A9", x"08", x"85", x"2C", x"38", x"20",
x"99", x"FF", x"C0", x"80", x"F0", x"03", x"A9", x"D0",
x"2C", x"A9", x"80", x"85", x"38", x"A9", x"00", x"85",
x"37", x"38", x"A5", x"37", x"E5", x"2B", x"AA", x"A5",
x"38", x"E5", x"2C", x"20", x"51", x"B4", x"A2", x"01",
x"4C", x"59", x"B9", x"05", x"05", x"06", x"06", x"08",
x"02", x"01", x"04", x"04", x"04", x"04", x"04", x"04",
x"07", x"03", x"C1", x"7B", x"53", x"F3", x"59", x"CC",
x"5C", x"74", x"35", x"AD", x"CF", x"AA", x"0E", x"BE",
x"BB", x"AA", x"BF", x"E4", x"BC", x"E0", x"BB", x"E0",
x"BF", x"BC", x"B1", x"BD", x"B1", x"E3", x"B8", x"B8",
x"EE", x"EF", x"F0", x"F1", x"F2", x"F3", x"F4", x"F5",
x"F6", x"F7", x"F8", x"F9", x"FA", x"FB", x"FC", x"FD",
x"FE", x"FF", x"00", x"01", x"02", x"03", x"04", x"E2",
x"E2", x"E2", x"E2", x"E2", x"E2", x"E2", x"E2", x"E2",
x"E2", x"E2", x"E2", x"E2", x"E2", x"E2", x"E2", x"E2",
x"E2", x"E3", x"E3", x"E3", x"E3", x"E3", x"08", x"18",
x"A5", x"2A", x"10", x"01", x"38", x"A5", x"29", x"85",
x"2A", x"A5", x"28", x"85", x"29", x"A5", x"27", x"85",
x"28", x"A5", x"26", x"85", x"27", x"A9", x"00", x"85",
x"26", x"90", x"12", x"E6", x"2A", x"D0", x"0E", x"E6",
x"29", x"D0", x"0A", x"E6", x"28", x"D0", x"06", x"E6",
x"27", x"D0", x"02", x"E6", x"26", x"28", x"60", x"84",
x"23", x"86", x"22", x"A0", x"00", x"A5", x"61", x"91",
x"22", x"F0", x"22", x"C8", x"A5", x"6D", x"91", x"22",
x"A5", x"66", x"D0", x"06", x"A5", x"6D", x"29", x"7F",
x"91", x"22", x"C8", x"A5", x"6C", x"91", x"22", x"C8",
x"A5", x"6B", x"91", x"22", x"C8", x"A5", x"6A", x"91",
x"22", x"A0", x"00", x"84", x"70", x"A5", x"61", x"60",
x"60", x"4C", x"B2", x"A6", x"20", x"4D", x"A1", x"38",
x"E9", x"AA", x"90", x"0E", x"C9", x"0A", x"B0", x"0A",
x"C9", x"07", x"F0", x"0B", x"C9", x"09", x"F0", x"19",
x"18", x"60", x"20", x"9C", x"A6", x"38", x"60", x"20",
x"4D", x"A1", x"C9", x"B2", x"F0", x"07", x"20", x"9C",
x"A6", x"A9", x"07", x"D0", x"EB", x"A9", x"0A", x"D0",
x"E7", x"20", x"4D", x"A1", x"C9", x"B2", x"F0", x"0B",
x"C9", x"B1", x"F0", x"0B", x"20", x"9C", x"A6", x"A9",
x"09", x"D0", x"D5", x"A9", x"0B", x"D0", x"D1", x"A9",
x"0C", x"D0", x"CD", x"60", x"38", x"A5", x"33", x"E5",
x"31", x"85", x"24", x"A5", x"34", x"E5", x"32", x"85",
x"25", x"90", x"1D", x"A5", x"24", x"E5", x"62", x"85",
x"24", x"A5", x"25", x"E5", x"63", x"85", x"25", x"90",
x"0F", x"A5", x"25", x"D0", x"0A", x"A5", x"61", x"0A",
x"18", x"69", x"04", x"C5", x"24", x"B0", x"01", x"60",
x"4C", x"CA", x"A6", x"60", x"A0", x"00", x"A2", x"5C",
x"4C", x"D4", x"BB", x"E6", x"61", x"D0", x"03", x"4C",
x"A3", x"B8", x"60", x"A5", x"91", x"30", x"03", x"4C",
x"90", x"A2", x"20", x"7F", x"AF", x"C9", x"3A", x"F0",
x"F9", x"C9", x"00", x"F0", x"44", x"AA", x"A9", x"A1",
x"48", x"A9", x"D9", x"48", x"E0", x"01", x"F0", x"1E",
x"E0", x"CB", x"D0", x"03", x"4C", x"8C", x"B4", x"E0",
x"7F", x"B0", x"03", x"4C", x"1F", x"A5", x"E0", x"A7",
x"90", x"03", x"4C", x"CF", x"A6", x"BD", x"26", x"BD",
x"48", x"BD", x"FF", x"BC", x"48", x"60", x"20", x"4D",
x"A1", x"C9", x"00", x"D0", x"03", x"4C", x"CF", x"A6",
x"C9", x"04", x"90", x"03", x"4C", x"CF", x"A6", x"AA",
x"BD", x"5E", x"B8", x"48", x"BD", x"5B", x"B8", x"48",
x"60", x"A6", x"3A", x"E8", x"D0", x"03", x"4C", x"34",
x"AC", x"A5", x"39", x"85", x"3B", x"A5", x"3A", x"85",
x"3C", x"20", x"32", x"E1", x"A5", x"3D", x"05", x"3E",
x"D0", x"03", x"4C", x"34", x"AC", x"20", x"A9", x"E3",
x"D0", x"03", x"4C", x"34", x"AC", x"A5", x"3D", x"18",
x"69", x"04", x"85", x"7A", x"A5", x"3E", x"69", x"00",
x"85", x"7B", x"A0", x"02", x"4C", x"80", x"E4", x"E0",
x"40", x"D0", x"03", x"4C", x"B8", x"A6", x"E0", x"5F",
x"D0", x"03", x"4C", x"B8", x"A6", x"20", x"9C", x"A6",
x"4C", x"F3", x"BD", x"20", x"12", x"BC", x"A0", x"01",
x"20", x"95", x"E1", x"C9", x"00", x"D0", x"01", x"60",
x"A0", x"04", x"20", x"95", x"E1", x"C9", x"00", x"F0",
x"06", x"C8", x"D0", x"F6", x"4C", x"C3", x"A6", x"C8",
x"98", x"18", x"65", x"3D", x"48", x"08", x"A0", x"00",
x"91", x"3D", x"28", x"A5", x"3E", x"69", x"00", x"A0",
x"01", x"91", x"3D", x"85", x"3E", x"68", x"85", x"3D",
x"4C", x"36", x"A5", x"A2", x"09", x"20", x"59", x"B9",
x"A2", x"08", x"AD", x"A6", x"02", x"F0", x"02", x"A2",
x"07", x"4C", x"59", x"B9", x"60", x"20", x"7F", x"AF",
x"C9", x"B2", x"F0", x"03", x"4C", x"CF", x"A6", x"60",
x"20", x"46", x"A7", x"90", x"01", x"60", x"24", x"0C",
x"10", x"03", x"4C", x"01", x"BD", x"20", x"AD", x"AE",
x"D0", x"03", x"4C", x"0D", x"B6", x"20", x"37", x"AB",
x"D0", x"03", x"4C", x"F6", x"BA", x"20", x"66", x"BF",
x"D0", x"03", x"4C", x"09", x"A4", x"A5", x"2D", x"85",
x"47", x"A5", x"2E", x"85", x"48", x"A5", x"48", x"C5",
x"30", x"D0", x"06", x"A5", x"47", x"C5", x"2F", x"F0",
x"14", x"20", x"39", x"E3", x"D0", x"07", x"A9", x"02",
x"20", x"D3", x"BD", x"18", x"60", x"A9", x"07", x"20",
x"D3", x"BD", x"4C", x"B5", x"A5", x"38", x"A5", x"33",
x"E5", x"31", x"48", x"A5", x"34", x"E5", x"32", x"D0",
x"08", x"68", x"C9", x"07", x"B0", x"04", x"4C", x"CA",
x"A6", x"68", x"38", x"A5", x"31", x"85", x"24", x"E5",
x"2F", x"85", x"28", x"A5", x"32", x"85", x"25", x"E5",
x"30", x"85", x"29", x"05", x"28", x"F0", x"16", x"E6",
x"28", x"D0", x"02", x"E6", x"29", x"18", x"A5", x"24",
x"69", x"07", x"85", x"26", x"A5", x"25", x"69", x"00",
x"85", x"27", x"20", x"A6", x"AD", x"18", x"A5", x"31",
x"69", x"07", x"85", x"31", x"90", x"02", x"E6", x"32",
x"18", x"A5", x"2F", x"69", x"07", x"85", x"2F", x"90",
x"02", x"E6", x"30", x"20", x"18", x"B4", x"A0", x"00",
x"A5", x"45", x"91", x"47", x"C8", x"A5", x"46", x"91",
x"47", x"C8", x"A9", x"00", x"91", x"47", x"C8", x"91",
x"47", x"4C", x"C6", x"A5", x"60", x"A9", x"25", x"20",
x"2E", x"BA", x"90", x"03", x"4C", x"CF", x"A6", x"A5",
x"15", x"C9", x"FF", x"D0", x"03", x"4C", x"B4", x"A6",
x"60", x"60", x"20", x"2E", x"BA", x"90", x"03", x"4C",
x"CF", x"A6", x"A5", x"14", x"48", x"A5", x"15", x"48",
x"20", x"C3", x"A1", x"90", x"03", x"4C", x"CF", x"A6",
x"48", x"20", x"C3", x"A1", x"90", x"02", x"A9", x"00",
x"85", x"25", x"68", x"85", x"24", x"68", x"85", x"23",
x"68", x"85", x"22", x"A0", x"00", x"B1", x"22", x"45",
x"25", x"25", x"24", x"F0", x"F8", x"60", x"A5", x"2B",
x"38", x"E9", x"01", x"85", x"7A", x"A5", x"2C", x"E9",
x"00", x"85", x"7B", x"60", x"A5", x"7A", x"38", x"E9",
x"01", x"85", x"7A", x"A5", x"7B", x"E9", x"00", x"85",
x"7B", x"60", x"AA", x"F0", x"0F", x"CA", x"10", x"3E",
x"E6", x"E6", x"E6", x"E6", x"E6", x"E6", x"E6", x"E6",
x"E6", x"E6", x"E6", x"E6", x"E6", x"E6", x"E6", x"E6",
x"E6", x"E6", x"E6", x"E6", x"E6", x"E6", x"E6", x"E6",
x"E6", x"E6", x"E6", x"E6", x"E6", x"E6", x"E6", x"E6",
x"E6", x"E6", x"E6", x"E6", x"E6", x"E6", x"E6", x"E6",
x"E6", x"EA", x"A5", x"E6", x"48", x"29", x"80", x"85",
x"E6", x"68", x"0A", x"05", x"EA", x"29", x"7F", x"AA",
x"A5", x"EA", x"29", x"80", x"85", x"EA", x"8A", x"48",
x"20", x"60", x"E0", x"A2", x"00", x"20", x"59", x"B9",
x"68", x"AA", x"20", x"53", x"B9", x"A2", x"03", x"20",
x"59", x"B9", x"A5", x"3A", x"C9", x"FF", x"F0", x"0C",
x"A2", x"04", x"20", x"59", x"B9", x"A5", x"3A", x"A6",
x"39", x"20", x"51", x"B4", x"A2", x"FE", x"9A", x"4C",
x"34", x"AC", x"60", x"20", x"7F", x"AF", x"C9", x"2C",
x"F0", x"05", x"20", x"9C", x"A6", x"38", x"60", x"18",
x"60", x"20", x"C1", x"B9", x"B0", x"17", x"20", x"AE",
x"AD", x"A5", x"0D", x"30", x"03", x"4C", x"CF", x"A6",
x"A5", x"61", x"85", x"B7", x"A5", x"62", x"85", x"BB",
x"A5", x"63", x"85", x"BC", x"18", x"60", x"A9", x"00",
x"85", x"46", x"20", x"7F", x"AF", x"20", x"76", x"A1",
x"90", x"05", x"20", x"9C", x"A6", x"38", x"60", x"85",
x"45", x"20", x"4D", x"A1", x"20", x"69", x"A1", x"B0",
x"0A", x"85", x"46", x"20", x"4D", x"A1", x"20", x"69",
x"A1", x"90", x"F8", x"C9", x"24", x"F0", x"1E", x"C9",
x"25", x"F0", x"0A", x"A9", x"05", x"85", x"53", x"20",
x"9C", x"A6", x"4C", x"9B", x"A7", x"A0", x"02", x"A9",
x"02", x"85", x"53", x"A5", x"45", x"09", x"80", x"85",
x"45", x"A9", x"00", x"F0", x"04", x"A0", x"03", x"A9",
x"FF", x"85", x"0D", x"84", x"53", x"A5", x"46", x"09",
x"80", x"85", x"46", x"20", x"7F", x"AF", x"C9", x"28",
x"F0", x"06", x"20", x"9C", x"A6", x"A9", x"00", x"2C",
x"A9", x"FF", x"85", x"0C", x"18", x"60", x"4C", x"96",
x"B4", x"A5", x"08", x"38", x"E5", x"07", x"18", x"69",
x"05", x"AA", x"20", x"57", x"E4", x"A0", x"01", x"98",
x"91", x"3D", x"C8", x"A5", x"14", x"91", x"3D", x"C8",
x"A5", x"15", x"91", x"3D", x"E6", x"08", x"A6", x"07",
x"BD", x"00", x"02", x"E6", x"07", x"C8", x"91", x"3D",
x"A5", x"07", x"C5", x"08", x"D0", x"F0", x"20", x"33",
x"A5", x"4C", x"12", x"E3", x"60", x"A0", x"0B", x"B9",
x"59", x"A1", x"99", x"00", x"03", x"88", x"10", x"F7",
x"A0", x"04", x"B9", x"65", x"A1", x"99", x"03", x"00",
x"88", x"10", x"F7", x"A9", x"4C", x"8D", x"10", x"03",
x"A9", x"CC", x"8D", x"11", x"03", x"A9", x"A6", x"8D",
x"12", x"03", x"A9", x"00", x"85", x"B0", x"85", x"B1",
x"20", x"22", x"E4", x"20", x"EB", x"B9", x"4C", x"B7",
x"E3", x"A5", x"62", x"C5", x"6A", x"90", x"3B", x"D0",
x"1D", x"A5", x"63", x"C5", x"6B", x"90", x"33", x"D0",
x"15", x"A5", x"64", x"C5", x"6C", x"90", x"2B", x"D0",
x"0D", x"A5", x"65", x"C5", x"6D", x"90", x"23", x"D0",
x"05", x"A9", x"00", x"85", x"61", x"60", x"38", x"A5",
x"65", x"E5", x"6D", x"85", x"65", x"A5", x"64", x"E5",
x"6C", x"85", x"64", x"A5", x"63", x"E5", x"6B", x"85",
x"63", x"A5", x"62", x"E5", x"6A", x"85", x"62", x"4C",
x"1E", x"B5", x"20", x"B8", x"BF", x"38", x"A9", x"00",
x"E5", x"70", x"85", x"70", x"A5", x"6D", x"E5", x"65",
x"85", x"65", x"A5", x"6C", x"E5", x"64", x"85", x"64",
x"A5", x"6B", x"E5", x"63", x"85", x"63", x"A5", x"6A",
x"E5", x"62", x"85", x"62", x"4C", x"1E", x"B5", x"A9",
x"00", x"9D", x"00", x"02", x"20", x"E7", x"FF", x"20",
x"59", x"F8", x"A9", x"0F", x"A0", x"0F", x"20", x"BA",
x"FF", x"20", x"45", x"BC", x"20", x"4D", x"A1", x"A0",
x"00", x"B1", x"7A", x"D0", x"03", x"4C", x"26", x"A9",
x"C9", x"24", x"D0", x"03", x"4C", x"45", x"A9", x"20",
x"6F", x"A1", x"90", x"23", x"20", x"B5", x"A9", x"20",
x"BD", x"FF", x"20", x"C0", x"FF", x"90", x"03", x"4C",
x"AD", x"A9", x"20", x"E7", x"FF", x"20", x"F1", x"A8",
x"AD", x"00", x"02", x"C9", x"30", x"D0", x"65", x"4D",
x"01", x"02", x"D0", x"60", x"4C", x"A7", x"A9", x"20",
x"C8", x"A1", x"C9", x"08", x"B0", x"03", x"4C", x"D1",
x"A6", x"48", x"20", x"7F", x"AF", x"C9", x"24", x"F0",
x"5F", x"C9", x"00", x"F0", x"03", x"4C", x"CF", x"A6",
x"68", x"85", x"BA", x"4C", x"34", x"AC", x"20", x"D2",
x"F7", x"A9", x"00", x"20", x"BD", x"FF", x"20", x"C0",
x"FF", x"90", x"03", x"4C", x"AD", x"A9", x"A2", x"0F",
x"20", x"C6", x"FF", x"90", x"03", x"4C", x"AD", x"A9",
x"A0", x"00", x"C0", x"50", x"D0", x"03", x"4C", x"CB",
x"A6", x"20", x"B7", x"FF", x"D0", x"0E", x"20", x"CF",
x"FF", x"90", x"03", x"4C", x"AD", x"A9", x"99", x"00",
x"02", x"C8", x"D0", x"E6", x"88", x"60", x"20", x"EE",
x"A8", x"4C", x"2F", x"A9", x"20", x"D2", x"F7", x"A2",
x"00", x"88", x"30", x"09", x"BD", x"00", x"02", x"20",
x"D2", x"FF", x"E8", x"D0", x"F4", x"4C", x"A7", x"A9",
x"68", x"85", x"BA", x"C6", x"7A", x"A9", x"00", x"A6",
x"BA", x"A0", x"60", x"20", x"BA", x"FF", x"20", x"B5",
x"A9", x"20", x"C0", x"FF", x"B0", x"57", x"A2", x"00",
x"20", x"C6", x"FF", x"B0", x"50", x"20", x"CF", x"FF",
x"B0", x"4B", x"20", x"CF", x"FF", x"B0", x"46", x"A0",
x"FF", x"C8", x"20", x"CF", x"FF", x"B0", x"3E", x"99",
x"00", x"02", x"C0", x"50", x"D0", x"03", x"4C", x"CB",
x"A6", x"20", x"B7", x"FF", x"D0", x"0B", x"C0", x"04",
x"90", x"E7", x"B9", x"00", x"02", x"D0", x"E2", x"F0",
x"04", x"A9", x"40", x"85", x"90", x"C0", x"05", x"90",
x"16", x"A9", x"00", x"99", x"00", x"02", x"A2", x"00",
x"86", x"3D", x"A2", x"02", x"86", x"3E", x"A2", x"3D",
x"20", x"85", x"AB", x"A5", x"90", x"F0", x"C0", x"20",
x"E7", x"FF", x"4C", x"34", x"AC", x"48", x"20", x"E7",
x"FF", x"68", x"4C", x"AA", x"A6", x"A0", x"FF", x"C8",
x"B1", x"7A", x"D0", x"FB", x"98", x"A6", x"7A", x"A4",
x"7B", x"4C", x"BD", x"FF", x"60", x"A9", x"00", x"85",
x"61", x"60", x"A5", x"61", x"F0", x"FB", x"A5", x"69",
x"D0", x"04", x"85", x"61", x"F0", x"F3", x"A5", x"66",
x"45", x"6E", x"85", x"66", x"20", x"95", x"A1", x"A5",
x"61", x"20", x"A2", x"A1", x"A5", x"69", x"20", x"A2",
x"A1", x"A5", x"26", x"E9", x"80", x"85", x"26", x"B0",
x"08", x"A5", x"27", x"E9", x"00", x"90", x"CE", x"85",
x"27", x"A5", x"27", x"F0", x"03", x"4C", x"A3", x"B8",
x"A5", x"26", x"85", x"61", x"20", x"95", x"A1", x"18",
x"A5", x"70", x"20", x"67", x"AA", x"20", x"A6", x"A3",
x"90", x"02", x"E6", x"26", x"A5", x"65", x"20", x"67",
x"AA", x"20", x"A6", x"A3", x"90", x"02", x"E6", x"26",
x"A5", x"64", x"20", x"67", x"AA", x"20", x"A6", x"A3",
x"90", x"02", x"E6", x"26", x"A5", x"63", x"20", x"67",
x"AA", x"20", x"A6", x"A3", x"90", x"02", x"E6", x"26",
x"A5", x"62", x"20", x"67", x"AA", x"20", x"A6", x"A3",
x"90", x"02", x"E6", x"26", x"A5", x"2A", x"85", x"70",
x"A5", x"29", x"85", x"65", x"A5", x"28", x"85", x"64",
x"A5", x"27", x"85", x"63", x"A5", x"26", x"85", x"62",
x"A5", x"61", x"18", x"69", x"08", x"90", x"03", x"4C",
x"A3", x"B8", x"85", x"61", x"4C", x"1E", x"B5", x"F0",
x"52", x"85", x"25", x"A5", x"6D", x"20", x"CD", x"BC",
x"65", x"2A", x"85", x"2A", x"8A", x"65", x"29", x"85",
x"29", x"90", x"0A", x"E6", x"28", x"D0", x"06", x"E6",
x"27", x"D0", x"02", x"E6", x"26", x"A5", x"6C", x"20",
x"CD", x"BC", x"65", x"29", x"85", x"29", x"8A", x"65",
x"28", x"85", x"28", x"90", x"06", x"E6", x"27", x"D0",
x"02", x"E6", x"26", x"A5", x"6B", x"20", x"CD", x"BC",
x"65", x"28", x"85", x"28", x"8A", x"65", x"27", x"85",
x"27", x"90", x"02", x"E6", x"26", x"A5", x"6A", x"20",
x"CD", x"BC", x"65", x"27", x"85", x"27", x"8A", x"65",
x"26", x"85", x"26", x"60", x"60", x"00", x"00", x"00",
x"03", x"27", x"68", x"45", x"0D", x"10", x"03", x"4C",
x"C4", x"A6", x"A5", x"0D", x"30", x"03", x"4C", x"B2",
x"A6", x"68", x"85", x"6B", x"68", x"85", x"6A", x"68",
x"85", x"69", x"F0", x"3C", x"A5", x"61", x"D0", x"12",
x"20", x"5C", x"BC", x"A5", x"69", x"85", x"61", x"A5",
x"6A", x"85", x"62", x"A5", x"6B", x"85", x"63", x"4C",
x"80", x"AE", x"18", x"65", x"69", x"90", x"03", x"4C",
x"C3", x"A6", x"20", x"07", x"E1", x"A0", x"01", x"B1",
x"47", x"85", x"22", x"C8", x"B1", x"47", x"85", x"23",
x"20", x"94", x"E4", x"20", x"5C", x"BC", x"A0", x"02",
x"B1", x"47", x"99", x"61", x"00", x"88", x"10", x"F8",
x"20", x"65", x"BC", x"4C", x"80", x"AE", x"84", x"36",
x"85", x"35", x"8A", x"48", x"A0", x"00", x"98", x"AA",
x"B1", x"35", x"F0", x"08", x"20", x"D2", x"FF", x"8A",
x"A8", x"C8", x"D0", x"F2", x"68", x"AA", x"60", x"A5",
x"46", x"C9", x"49", x"D0", x"04", x"A5", x"45", x"C9",
x"54", x"60", x"A2", x"20", x"06", x"6D", x"26", x"6C",
x"26", x"6B", x"26", x"6A", x"26", x"29", x"26", x"28",
x"26", x"27", x"26", x"26", x"38", x"A5", x"29", x"E5",
x"65", x"85", x"25", x"A5", x"28", x"E5", x"64", x"85",
x"24", x"A5", x"27", x"E5", x"63", x"85", x"23", x"A5",
x"26", x"E5", x"62", x"90", x"14", x"85", x"22", x"A5",
x"25", x"85", x"29", x"A5", x"24", x"85", x"28", x"A5",
x"23", x"85", x"27", x"A5", x"22", x"85", x"26", x"E6",
x"6D", x"CA", x"D0", x"C0", x"60", x"20", x"D2", x"F7",
x"A0", x"03", x"20", x"95", x"E1", x"48", x"88", x"20",
x"95", x"E1", x"AA", x"68", x"20", x"51", x"B4", x"20",
x"D7", x"F7", x"A9", x"00", x"85", x"D4", x"A0", x"04",
x"20", x"95", x"E1", x"C9", x"00", x"D0", x"01", x"60",
x"C9", x"22", x"D0", x"0B", x"A5", x"D4", x"49", x"FF",
x"85", x"D4", x"A9", x"22", x"4C", x"E4", x"AB", x"A6",
x"D4", x"D0", x"29", x"C9", x"FF", x"F0", x"23", x"C9",
x"01", x"F0", x"4F", x"C9", x"7F", x"90", x"1D", x"AA",
x"48", x"98", x"48", x"8A", x"29", x"7F", x"AA", x"E0",
x"4C", x"B0", x"3A", x"20", x"65", x"B9", x"68", x"A8",
x"68", x"C9", x"8F", x"D0", x"02", x"85", x"D4", x"C8",
x"D0", x"BE", x"A9", x"7E", x"48", x"24", x"D4", x"10",
x"19", x"29", x"7F", x"C9", x"12", x"F0", x"13", x"29",
x"60", x"D0", x"0F", x"68", x"98", x"48", x"A9", x"88",
x"A0", x"AF", x"20", x"1E", x"AB", x"68", x"A8", x"4C",
x"06", x"AC", x"68", x"20", x"D2", x"FF", x"C8", x"F0",
x"03", x"4C", x"A0", x"AB", x"60", x"68", x"68", x"4C",
x"F4", x"AB", x"20", x"23", x"AC", x"E0", x"03", x"B0",
x"DB", x"98", x"48", x"20", x"5F", x"B9", x"68", x"A8",
x"4C", x"DF", x"AB", x"C8", x"20", x"95", x"E1", x"C9",
x"00", x"AA", x"F0", x"02", x"CA", x"60", x"88", x"4C",
x"0D", x"AC", x"48", x"48", x"A2", x"02", x"20", x"59",
x"B9", x"A9", x"FF", x"85", x"3A", x"A9", x"80", x"20",
x"90", x"FF", x"A2", x"00", x"20", x"CF", x"FF", x"B0",
x"FB", x"C9", x"0D", x"F0", x"0E", x"E0", x"50", x"90",
x"03", x"4C", x"C3", x"A6", x"9D", x"00", x"02", x"E8",
x"4C", x"44", x"AC", x"86", x"07", x"A9", x"00", x"9D",
x"00", x"02", x"AD", x"00", x"02", x"C9", x"20", x"D0",
x"11", x"A2", x"01", x"BD", x"00", x"02", x"9D", x"FF",
x"01", x"E8", x"E4", x"07", x"D0", x"F5", x"C6", x"07",
x"D0", x"E8", x"20", x"D2", x"F7", x"A5", x"07", x"F0",
x"C1", x"A6", x"07", x"AD", x"00", x"02", x"C9", x"40",
x"D0", x"03", x"4C", x"7F", x"A8", x"C9", x"5F", x"D0",
x"03", x"4C", x"7F", x"A1", x"20", x"62", x"B6", x"AD",
x"00", x"02", x"C9", x"30", x"90", x"43", x"C9", x"3A",
x"B0", x"3F", x"A5", x"07", x"85", x"08", x"A9", x"00",
x"85", x"07", x"A9", x"00", x"85", x"7A", x"A9", x"02",
x"85", x"7B", x"20", x"45", x"A6", x"A5", x"7A", x"85",
x"07", x"A6", x"07", x"BD", x"00", x"02", x"C9", x"20",
x"D0", x"03", x"E8", x"D0", x"F6", x"86", x"07", x"20",
x"12", x"E3", x"20", x"14", x"E2", x"B0", x"06", x"20",
x"F1", x"A2", x"20", x"14", x"E2", x"A5", x"07", x"C5",
x"08", x"F0", x"03", x"20", x"B1", x"A7", x"4C", x"42",
x"AC", x"20", x"45", x"BC", x"4C", x"93", x"A4", x"A9",
x"00", x"A0", x"1D", x"99", x"01", x"01", x"88", x"10",
x"FA", x"BD", x"00", x"02", x"C9", x"23", x"90", x"20",
x"C9", x"7B", x"B0", x"1C", x"C9", x"30", x"90", x"04",
x"C9", x"3C", x"90", x"14", x"A0", x"0E", x"D9", x"B0",
x"B1", x"F0", x"0E", x"88", x"D0", x"F8", x"A0", x"16",
x"D9", x"57", x"A2", x"F0", x"43", x"88", x"D0", x"F8",
x"60", x"2C", x"04", x"01", x"10", x"2E", x"98", x"0A",
x"0A", x"0A", x"0A", x"AC", x"05", x"01", x"19", x"06",
x"01", x"99", x"06", x"01", x"EE", x"05", x"01", x"EE",
x"04", x"01", x"18", x"6E", x"02", x"01", x"6E", x"03",
x"01", x"E8", x"EE", x"01", x"01", x"AD", x"01", x"01",
x"C9", x"07", x"F0", x"07", x"BD", x"FF", x"01", x"C9",
x"41", x"B0", x"A6", x"60", x"98", x"AC", x"05", x"01",
x"99", x"06", x"01", x"CE", x"04", x"01", x"30", x"DA",
x"2C", x"04", x"01", x"10", x"22", x"98", x"48", x"A9",
x"F0", x"AC", x"05", x"01", x"19", x"06", x"01", x"99",
x"06", x"01", x"C8", x"68", x"99", x"06", x"01", x"C8",
x"8C", x"05", x"01", x"EE", x"04", x"01", x"38", x"6E",
x"02", x"01", x"6E", x"03", x"01", x"90", x"BA", x"98",
x"AC", x"05", x"01", x"99", x"06", x"01", x"C8", x"29",
x"0F", x"99", x"06", x"01", x"88", x"B9", x"06", x"01",
x"09", x"0F", x"99", x"06", x"01", x"C8", x"8C", x"05",
x"01", x"CE", x"04", x"01", x"30", x"D8", x"4C", x"AE",
x"AD", x"01", x"0A", x"64", x"E8", x"10", x"A4", x"28",
x"20", x"3D", x"A2", x"4C", x"B0", x"E1", x"A9", x"00",
x"48", x"20", x"C1", x"B9", x"90", x"03", x"4C", x"CF",
x"A6", x"20", x"4D", x"A1", x"C9", x"22", x"F0", x"56",
x"C9", x"28", x"F0", x"32", x"C9", x"AB", x"D0", x"03",
x"4C", x"F1", x"AD", x"C9", x"A8", x"D0", x"03", x"4C",
x"EE", x"AD", x"C9", x"FF", x"D0", x"03", x"4C", x"03",
x"AE", x"C9", x"80", x"B0", x"0E", x"20", x"9C", x"A6",
x"20", x"88", x"A5", x"B0", x"28", x"20", x"4D", x"E3",
x"4C", x"3A", x"AE", x"4C", x"B2", x"A6", x"A0", x"0D",
x"2C", x"A0", x"0E", x"4C", x"6A", x"AE", x"20", x"AE",
x"AD", x"20", x"4D", x"A1", x"C9", x"29", x"F0", x"3A",
x"4C", x"CF", x"A6", x"A9", x"A8", x"A0", x"AE", x"20",
x"9C", x"BC", x"4C", x"10", x"AE", x"4C", x"B2", x"A6",
x"A9", x"00", x"85", x"0D", x"F0", x"24", x"A2", x"FF",
x"86", x"0D", x"E8", x"86", x"61", x"A6", x"7A", x"86",
x"62", x"A6", x"7B", x"86", x"63", x"20", x"4D", x"A1",
x"C9", x"22", x"F0", x"0E", x"C9", x"00", x"F0", x"07",
x"E6", x"61", x"D0", x"F1", x"4C", x"C3", x"A6", x"20",
x"9C", x"A6", x"20", x"C1", x"B9", x"B0", x"3D", x"20",
x"0C", x"A4", x"B0", x"38", x"A8", x"68", x"48", x"D9",
x"4B", x"A3", x"90", x"0F", x"84", x"4C", x"A9", x"FF",
x"85", x"4B", x"4C", x"84", x"AE", x"68", x"48", x"D0",
x"F9", x"A4", x"4C", x"A6", x"0D", x"30", x"00", x"A5",
x"61", x"48", x"A5", x"62", x"48", x"A5", x"63", x"48",
x"8A", x"48", x"20", x"1E", x"BC", x"B9", x"69", x"A3",
x"48", x"B9", x"5A", x"A3", x"48", x"B9", x"4B", x"A3",
x"48", x"4C", x"B1", x"AD", x"A9", x"00", x"85", x"4B",
x"A5", x"4B", x"D0", x"D1", x"68", x"60", x"60", x"A5",
x"61", x"85", x"69", x"F0", x"16", x"A5", x"62", x"85",
x"6A", x"A5", x"63", x"85", x"6B", x"A5", x"64", x"85",
x"6C", x"A5", x"65", x"85", x"6D", x"A5", x"66", x"85",
x"6E", x"A5", x"61", x"A2", x"00", x"86", x"70", x"60",
x"82", x"49", x"0F", x"DA", x"A2", x"A5", x"46", x"C9",
x"C9", x"D0", x"04", x"A5", x"45", x"C9", x"54", x"60",
x"20", x"46", x"A7", x"90", x"03", x"4C", x"CF", x"A6",
x"20", x"95", x"B7", x"B0", x"03", x"4C", x"C7", x"A6",
x"A5", x"46", x"48", x"A5", x"45", x"48", x"A5", x"53",
x"48", x"24", x"0C", x"30", x"0A", x"A9", x"0A", x"48",
x"A9", x"00", x"48", x"A2", x"01", x"D0", x"1B", x"A2",
x"00", x"E8", x"20", x"74", x"A2", x"E6", x"14", x"D0",
x"02", x"E6", x"15", x"D0", x"03", x"4C", x"CA", x"A6",
x"A5", x"14", x"48", x"A5", x"15", x"48", x"C0", x"00",
x"F0", x"E7", x"8A", x"48", x"20", x"A3", x"AF", x"A0",
x"01", x"84", x"62", x"88", x"84", x"63", x"68", x"85",
x"61", x"20", x"54", x"A4", x"A5", x"61", x"A0", x"04",
x"91", x"31", x"C8", x"AA", x"68", x"91", x"31", x"85",
x"65", x"C8", x"68", x"91", x"31", x"85", x"64", x"C8",
x"20", x"01", x"B9", x"CA", x"D0", x"EE", x"84", x"66",
x"68", x"85", x"53", x"85", x"64", x"86", x"65", x"20",
x"01", x"B9", x"20", x"54", x"A4", x"A0", x"00", x"68",
x"91", x"31", x"C8", x"68", x"91", x"31", x"A9", x"05",
x"20", x"89", x"E0", x"A5", x"61", x"0A", x"20", x"89",
x"E0", x"A0", x"02", x"A5", x"22", x"91", x"31", x"C8",
x"A5", x"23", x"91", x"31", x"18", x"A5", x"66", x"65",
x"31", x"85", x"31", x"90", x"02", x"E6", x"32", x"A0",
x"00", x"A9", x"00", x"91", x"31", x"E6", x"31", x"D0",
x"02", x"E6", x"32", x"38", x"A5", x"62", x"E9", x"01",
x"85", x"62", x"B0", x"02", x"C6", x"63", x"05", x"63",
x"D0", x"E7", x"60", x"60", x"00", x"00", x"60", x"20",
x"4D", x"A1", x"C9", x"20", x"F0", x"F9", x"60", x"60",
x"12", x"3F", x"92", x"00", x"85", x"50", x"38", x"A5",
x"7A", x"E5", x"50", x"85", x"7A", x"B0", x"02", x"C6",
x"7B", x"60", x"60", x"20", x"C3", x"A1", x"B0", x"02",
x"85", x"B9", x"60", x"A5", x"7A", x"48", x"A5", x"7B",
x"48", x"A5", x"3D", x"48", x"A5", x"3E", x"48", x"A9",
x"00", x"85", x"22", x"85", x"23", x"A5", x"37", x"85",
x"7A", x"A5", x"38", x"85", x"7B", x"A5", x"34", x"C5",
x"7B", x"D0", x"20", x"A5", x"33", x"C5", x"7A", x"D0",
x"1A", x"18", x"A5", x"22", x"65", x"33", x"85", x"33",
x"A5", x"23", x"65", x"34", x"85", x"34", x"68", x"85",
x"3E", x"68", x"85", x"3D", x"68", x"85", x"7B", x"68",
x"85", x"7A", x"60", x"A9", x"02", x"20", x"8C", x"AF",
x"20", x"2F", x"E0", x"D0", x"03", x"4C", x"70", x"B0",
x"A0", x"00", x"20", x"95", x"E1", x"85", x"28", x"A9",
x"00", x"85", x"29", x"18", x"A5", x"28", x"69", x"02",
x"85", x"28", x"90", x"02", x"E6", x"29", x"C8", x"20",
x"66", x"E3", x"18", x"A5", x"24", x"65", x"28", x"85",
x"24", x"A5", x"25", x"65", x"29", x"85", x"25", x"38",
x"A5", x"24", x"E9", x"01", x"85", x"24", x"B0", x"02",
x"C6", x"25", x"18", x"A5", x"24", x"65", x"22", x"85",
x"26", x"A5", x"25", x"65", x"23", x"85", x"27", x"A0",
x"01", x"20", x"76", x"E3", x"20", x"A6", x"AD", x"A0",
x"00", x"20", x"95", x"E1", x"20", x"8C", x"AF", x"A5",
x"63", x"C5", x"7B", x"D0", x"11", x"A5", x"62", x"C5",
x"7A", x"D0", x"0B", x"18", x"65", x"22", x"85", x"62",
x"A5", x"63", x"65", x"23", x"85", x"63", x"A5", x"6B",
x"C5", x"7B", x"D0", x"11", x"A5", x"6A", x"C5", x"7A",
x"D0", x"0B", x"18", x"65", x"22", x"85", x"6A", x"A5",
x"6B", x"65", x"23", x"85", x"6B", x"4C", x"BD", x"AF",
x"A9", x"01", x"20", x"8C", x"AF", x"A0", x"00", x"20",
x"88", x"E1", x"AA", x"A9", x"03", x"20", x"89", x"E0",
x"8A", x"20", x"89", x"E0", x"8A", x"20", x"8C", x"AF",
x"4C", x"BD", x"AF", x"CD", x"05", x"00", x"A3", x"09",
x"00", x"DC", x"0F", x"ED", x"00", x"85", x"8E", x"00",
x"C7", x"26", x"FE", x"0A", x"00", x"C7", x"26", x"0E",
x"00", x"75", x"1F", x"03", x"00", x"D9", x"58", x"00",
x"D4", x"0E", x"00", x"1F", x"A5", x"AE", x"00", x"29",
x"0C", x"00", x"37", x"00", x"D9", x"EB", x"9A", x"0D",
x"00", x"1F", x"A5", x"2B", x"1F", x"02", x"00", x"D9",
x"2E", x"C9", x"00", x"D9", x"1F", x"03", x"00", x"EB",
x"6A", x"00", x"CA", x"00", x"0F", x"8F", x"E7", x"00",
x"A4", x"58", x"00", x"8B", x"1F", x"D1", x"00", x"1F",
x"D1", x"79", x"F3", x"0E", x"00", x"D5", x"03", x"00",
x"A6", x"0F", x"DC", x"00", x"96", x"C7", x"FE", x"0A",
x"00", x"96", x"C7", x"0E", x"00", x"1F", x"A6", x"EC",
x"00", x"74", x"EB", x"00", x"1F", x"46", x"09", x"00",
x"1F", x"F6", x"13", x"05", x"00", x"FB", x"0E", x"0B",
x"00", x"6A", x"CD", x"00", x"1F", x"46", x"BA", x"0D",
x"00", x"1F", x"D5", x"0E", x"00", x"DC", x"0F", x"0F",
x"00", x"8E", x"1F", x"F2", x"0B", x"00", x"AE", x"00",
x"C3", x"00", x"6B", x"1F", x"F6", x"0B", x"00", x"FE",
x"10", x"CD", x"00", x"AC", x"0E", x"00", x"EB", x"6D",
x"00", x"0F", x"08", x"00", x"0F", x"05", x"00", x"0F",
x"06", x"00", x"0F", x"04", x"00", x"0F", x"07", x"00",
x"C8", x"05", x"00", x"9A", x"00", x"0F", x"01", x"00",
x"0F", x"02", x"00", x"0F", x"03", x"00", x"FB", x"15",
x"0C", x"00", x"C7", x"0E", x"00", x"F8", x"12", x"0B",
x"00", x"B2", x"09", x"00", x"93", x"0D", x"00", x"A6",
x"0B", x"00", x"FB", x"09", x"09", x"00", x"C9", x"05",
x"00", x"A4", x"1F", x"05", x"00", x"FD", x"0D", x"06",
x"00", x"1F", x"A6", x"0B", x"00", x"7B", x"0C", x"00",
x"8E", x"0C", x"00", x"E8", x"0C", x"00", x"D6", x"FD",
x"0C", x"00", x"D4", x"0C", x"00", x"EB", x"F9", x"14",
x"00", x"1F", x"81", x"04", x"00", x"B8", x"1F", x"06",
x"00", x"1F", x"F6", x"10", x"F9", x"14", x"00", x"D4",
x"E3", x"1F", x"04", x"00", x"79", x"1F", x"F5", x"10",
x"FE", x"14", x"00", x"1F", x"73", x"F5", x"14", x"00",
x"1F", x"A5", x"00", x"FF", x"FF", x"90", x"80", x"00",
x"00", x"00", x"60", x"4C", x"B2", x"A6", x"4C", x"B2",
x"A6", x"20", x"55", x"46", x"4C", x"44", x"50", x"49",
x"41", x"52", x"4F", x"53", x"4E", x"45", x"54", x"60",
x"A6", x"3A", x"E8", x"F0", x"03", x"4C", x"B8", x"A6",
x"A0", x"01", x"98", x"91", x"2B", x"20", x"DE", x"A7",
x"4C", x"32", x"AC", x"1F", x"F7", x"1C", x"00", x"F1",
x"12", x"B8", x"F7", x"16", x"F1", x"12", x"0F", x"EE",
x"BD", x"31", x"D9", x"0D", x"00", x"1F", x"97", x"8D",
x"F5", x"0E", x"1F", x"FA", x"17", x"00", x"D1", x"99",
x"9A", x"00", x"71", x"1C", x"00", x"00", x"1F", x"F7",
x"12", x"F9", x"0C", x"81", x"1E", x"1F", x"04", x"00",
x"86", x"F4", x"17", x"00", x"EC", x"FB", x"16", x"1F",
x"07", x"00", x"8E", x"D6", x"41", x"8A", x"15", x"AC",
x"F9", x"13", x"48", x"E1", x"92", x"1F", x"A2", x"1F",
x"77", x"FD", x"16", x"51", x"4A", x"F6", x"10", x"C7",
x"F1", x"1B", x"37", x"F3", x"0E", x"1F", x"07", x"00",
x"D9", x"D4", x"B8", x"1D", x"00", x"AE", x"1A", x"1F",
x"83", x"FC", x"0E", x"31", x"47", x"BD", x"00", x"73",
x"D4", x"A1", x"D6", x"0C", x"00", x"73", x"D4", x"C1",
x"EA", x"A1", x"D6", x"0C", x"00", x"73", x"D4", x"C1",
x"EA", x"31", x"2A", x"5C", x"00", x"D5", x"1F", x"71",
x"1F", x"D6", x"C1", x"EA", x"61", x"D9", x"DB", x"EC",
x"00", x"AC", x"1E", x"C7", x"26", x"1E", x"73", x"D4",
x"00", x"AC", x"1E", x"2A", x"6E", x"E2", x"31", x"47",
x"0D", x"00", x"1F", x"73", x"BB", x"C7", x"1F", x"15",
x"73", x"D4", x"8C", x"1F", x"D3", x"00", x"47", x"D4",
x"1F", x"85", x"14", x"D5", x"1F", x"71", x"1F", x"D6",
x"C1", x"F2", x"13", x"1F", x"D2", x"09", x"00", x"DC",
x"0F", x"ED", x"F1", x"0F", x"E7", x"1F", x"A0", x"E2",
x"31", x"9A", x"00", x"FB", x"0E", x"EC", x"F8", x"0D",
x"00", x"D9", x"2E", x"C9", x"F1", x"0F", x"E7", x"1F",
x"A0", x"E2", x"F1", x"15", x"BA", x"F2", x"12", x"00",
x"2A", x"1E", x"3A", x"51", x"E8", x"08", x"00", x"47",
x"D4", x"1F", x"85", x"14", x"0F", x"29", x"C8", x"7E",
x"FE", x"0E", x"00", x"FA", x"11", x"9D", x"43", x"FA",
x"0F", x"00", x"2A", x"1E", x"3A", x"F1", x"13", x"FD",
x"13", x"9A", x"0F", x"0E", x"00", x"C2", x"D5", x"F3",
x"18", x"15", x"EB", x"E8", x"FD", x"13", x"CD", x"0E",
x"00", x"1F", x"82", x"15", x"2B", x"1F", x"B2", x"1F",
x"96", x"67", x"0E", x"00", x"D9", x"75", x"1F", x"F3",
x"18", x"15", x"98", x"89", x"0F", x"0E", x"00", x"75",
x"1F", x"71", x"7B", x"CA", x"F1", x"12", x"0F", x"1E",
x"1F", x"D9", x"A9", x"00", x"47", x"D4", x"1F", x"85",
x"14", x"75", x"D9", x"1F", x"E6", x"00", x"FE", x"0E",
x"D6", x"F1", x"13", x"B7", x"1F", x"83", x"FE", x"16",
x"1F", x"00", x"EB", x"79", x"FC", x"15", x"E1", x"AA",
x"41", x"CA", x"1F", x"05", x"00", x"73", x"D4", x"51",
x"E8", x"08", x"00", x"A3", x"F9", x"13", x"42", x"18",
x"AE", x"1A", x"1F", x"A6", x"1F", x"63", x"D4", x"0F",
x"0D", x"00", x"1F", x"86", x"FC", x"18", x"1E", x"1F",
x"A6", x"EC", x"C7", x"D2", x"00", x"C2", x"D5", x"F3",
x"18", x"15", x"23", x"FC", x"16", x"7E", x"CA", x"00",
x"1F", x"D1", x"79", x"F3", x"0E", x"00", x"A4", x"58",
x"00", x"1F", x"92", x"8D", x"0F", x"0C", x"00", x"00",
x"00", x"00", x"75", x"D9", x"1F", x"E6", x"F1", x"13",
x"5A", x"1D", x"CA", x"F4", x"0E", x"00", x"00", x"00",
x"00", x"74", x"DC", x"C1", x"F2", x"13", x"1F", x"D2",
x"19", x"AE", x"1A", x"84", x"F9", x"15", x"0D", x"00",
x"00", x"AC", x"1E", x"F7", x"13", x"46", x"FD", x"13",
x"CD", x"DE", x"05", x"00", x"00", x"1F", x"D3", x"1F",
x"A3", x"F9", x"0E", x"F1", x"16", x"9A", x"29", x"E6",
x"00", x"60", x"8D", x"7A", x"D0", x"A9", x"00", x"F0",
x"05", x"8D", x"7B", x"D0", x"A9", x"01", x"8D", x"30",
x"D0", x"60", x"60", x"18", x"A5", x"33", x"65", x"50",
x"85", x"33", x"90", x"02", x"E6", x"34", x"60", x"A5",
x"50", x"D0", x"01", x"60", x"20", x"48", x"B9", x"B0",
x"01", x"60", x"D0", x"0A", x"20", x"A3", x"B3", x"A9",
x"02", x"85", x"50", x"4C", x"A3", x"B3", x"C6", x"50",
x"18", x"A5", x"51", x"65", x"50", x"85", x"51", x"90",
x"02", x"E6", x"52", x"A5", x"50", x"A0", x"00", x"91",
x"51", x"98", x"C8", x"91", x"51", x"C8", x"91", x"51",
x"60", x"20", x"7F", x"AF", x"C9", x"00", x"F0", x"25",
x"C9", x"22", x"F0", x"03", x"4C", x"CF", x"A6", x"A5",
x"7A", x"85", x"BB", x"A5", x"7B", x"85", x"BC", x"A2",
x"00", x"20", x"4D", x"A1", x"C9", x"00", x"F0", x"07",
x"C9", x"22", x"F0", x"03", x"E8", x"D0", x"F2", x"86",
x"B7", x"A9", x"00", x"F0", x"02", x"85", x"B7", x"85",
x"0A", x"A0", x"01", x"A2", x"07", x"4C", x"BA", x"FF",
x"A5", x"2F", x"85", x"22", x"A5", x"30", x"85", x"23",
x"A5", x"23", x"C5", x"32", x"D0", x"07", x"A5", x"22",
x"C5", x"31", x"D0", x"01", x"60", x"20", x"E1", x"E1",
x"B0", x"14", x"20", x"63", x"E1", x"A9", x"03", x"20",
x"89", x"E0", x"A5", x"22", x"C5", x"24", x"D0", x"F2",
x"A5", x"23", x"C5", x"25", x"D0", x"EC", x"A5", x"25",
x"85", x"23", x"A5", x"24", x"85", x"22", x"4C", x"20",
x"B4", x"85", x"62", x"86", x"61", x"05", x"61", x"D0",
x"05", x"A9", x"30", x"4C", x"D2", x"FF", x"A0", x"04",
x"20", x"FF", x"BB", x"B0", x"03", x"88", x"10", x"F8",
x"A2", x"00", x"20", x"FF", x"BB", x"90", x"12", x"E8",
x"38", x"A5", x"61", x"F9", x"A1", x"AD", x"85", x"61",
x"A5", x"62", x"F9", x"BD", x"AA", x"85", x"62", x"B0",
x"E9", x"8A", x"18", x"69", x"30", x"20", x"D2", x"FF",
x"88", x"10", x"DD", x"60", x"20", x"7F", x"AF", x"C9",
x"A4", x"F0", x"13", x"4C", x"CF", x"A6", x"20", x"00",
x"BA", x"20", x"12", x"BC", x"A9", x"00", x"20", x"90",
x"FF", x"20", x"C1", x"B9", x"B0", x"28", x"20", x"45",
x"A6", x"B0", x"E8", x"A5", x"3A", x"30", x"12", x"A5",
x"15", x"C5", x"3A", x"D0", x"04", x"A5", x"14", x"C5",
x"39", x"90", x"0B", x"20", x"17", x"E2", x"4C", x"C9",
x"B4", x"A9", x"00", x"20", x"90", x"FF", x"20", x"14",
x"E2", x"90", x"03", x"4C", x"C9", x"A6", x"48", x"48",
x"4C", x"05", x"A5", x"A9", x"00", x"85", x"0F", x"A5",
x"33", x"85", x"22", x"A5", x"34", x"85", x"23", x"A9",
x"02", x"20", x"09", x"A2", x"B0", x"21", x"A0", x"00",
x"A5", x"47", x"91", x"33", x"C8", x"A5", x"48", x"91",
x"33", x"A0", x"00", x"20", x"9E", x"E1", x"20", x"09",
x"A2", x"B0", x"0C", x"A0", x"01", x"A5", x"33", x"91",
x"47", x"C8", x"A5", x"34", x"91", x"47", x"60", x"A5",
x"22", x"85", x"33", x"A5", x"23", x"85", x"34", x"24",
x"0F", x"30", x"03", x"4C", x"CA", x"A6", x"C6", x"0F",
x"20", x"A3", x"AF", x"4C", x"D5", x"B4", x"A5", x"61",
x"F0", x"48", x"A5", x"62", x"F0", x"17", x"A5", x"62",
x"29", x"80", x"D0", x"3E", x"C6", x"61", x"F0", x"3A",
x"06", x"70", x"26", x"65", x"26", x"64", x"26", x"63",
x"26", x"62", x"90", x"EA", x"60", x"A5", x"61", x"38",
x"E9", x"08", x"B0", x"02", x"A9", x"00", x"85", x"61",
x"F0", x"20", x"A5", x"63", x"85", x"62", x"A5", x"64",
x"85", x"63", x"A5", x"65", x"85", x"64", x"A5", x"70",
x"85", x"65", x"A9", x"00", x"85", x"70", x"05", x"62",
x"05", x"63", x"05", x"64", x"05", x"65", x"D0", x"BA",
x"85", x"61", x"60", x"CE", x"01", x"01", x"F0", x"1F",
x"0E", x"03", x"01", x"2E", x"02", x"01", x"B0", x"21",
x"AC", x"05", x"01", x"2C", x"04", x"01", x"30", x"10",
x"88", x"8C", x"05", x"01", x"B9", x"06", x"01", x"29",
x"0F", x"99", x"06", x"01", x"CE", x"04", x"01", x"60",
x"A9", x"00", x"99", x"06", x"01", x"EE", x"04", x"01",
x"60", x"AC", x"05", x"01", x"A9", x"00", x"2C", x"04",
x"01", x"30", x"0A", x"88", x"99", x"06", x"01", x"8C",
x"05", x"01", x"4C", x"80", x"B5", x"99", x"06", x"01",
x"88", x"99", x"06", x"01", x"8C", x"05", x"01", x"EE",
x"04", x"01", x"60", x"20", x"C1", x"B9", x"90", x"03",
x"4C", x"CF", x"A6", x"A0", x"00", x"B1", x"7A", x"D9",
x"07", x"B6", x"D0", x"11", x"B1", x"7A", x"F0", x"03",
x"C8", x"D0", x"F2", x"A9", x"0C", x"85", x"14", x"A9",
x"08", x"85", x"15", x"D0", x"0A", x"A9", x"0A", x"20",
x"2E", x"BA", x"90", x"03", x"4C", x"CF", x"A6", x"A9",
x"4C", x"8D", x"10", x"03", x"A5", x"14", x"8D", x"11",
x"03", x"A5", x"15", x"8D", x"12", x"03", x"AD", x"0F",
x"03", x"48", x"AC", x"0E", x"03", x"AE", x"0D", x"03",
x"AD", x"0C", x"03", x"28", x"4C", x"10", x"03", x"FF",
x"AC", x"36", x"35", x"36", x"00", x"A9", x"06", x"20",
x"07", x"E1", x"20", x"EB", x"E3", x"20", x"DE", x"FF",
x"84", x"24", x"86", x"23", x"85", x"22", x"A0", x"00",
x"A9", x"30", x"85", x"25", x"A5", x"24", x"D9", x"CD",
x"E4", x"90", x"2C", x"D0", x"10", x"A5", x"23", x"D9",
x"09", x"BB", x"90", x"23", x"D0", x"07", x"A5", x"22",
x"D9", x"65", x"E2", x"90", x"1A", x"E6", x"25", x"38",
x"A5", x"22", x"F9", x"65", x"E2", x"85", x"22", x"A5",
x"23", x"F9", x"09", x"BB", x"85", x"23", x"A5", x"24",
x"F9", x"CD", x"E4", x"85", x"24", x"B0", x"CD", x"A5",
x"25", x"91", x"51", x"C8", x"C0", x"06", x"D0", x"C0",
x"18", x"60", x"A9", x"00", x"8D", x"00", x"01", x"A6",
x"07", x"9D", x"00", x"02", x"AD", x"00", x"01", x"C5",
x"07", x"F0", x"4D", x"AE", x"00", x"01", x"BD", x"00",
x"02", x"C9", x"22", x"F0", x"44", x"C9", x"DE", x"F0",
x"51", x"C9", x"3F", x"F0", x"50", x"20", x"E7", x"AC",
x"AD", x"01", x"01", x"F0", x"4D", x"A9", x"8B", x"85",
x"35", x"A9", x"B0", x"85", x"36", x"20", x"65", x"BB",
x"90", x"13", x"A9", x"C0", x"85", x"35", x"A9", x"E3",
x"85", x"36", x"20", x"65", x"BB", x"90", x"39", x"20",
x"6B", x"B5", x"4C", x"88", x"B6", x"8A", x"48", x"AE",
x"00", x"01", x"18", x"69", x"80", x"9D", x"00", x"02",
x"20", x"8E", x"E2", x"68", x"C9", x"0F", x"D0", x"AC",
x"60", x"EE", x"00", x"01", x"AE", x"00", x"01", x"BD",
x"00", x"02", x"F0", x"F4", x"C9", x"22", x"F0", x"0A",
x"D0", x"EF", x"A9", x"FF", x"2C", x"A9", x"99", x"9D",
x"00", x"02", x"EE", x"00", x"01", x"4C", x"6C", x"B6",
x"A9", x"01", x"AC", x"00", x"01", x"99", x"00", x"02",
x"E8", x"8A", x"C8", x"8C", x"00", x"01", x"99", x"00",
x"02", x"20", x"8B", x"E2", x"4C", x"6C", x"B6", x"A5",
x"61", x"C5", x"69", x"F0", x"50", x"B0", x"4F", x"A5",
x"69", x"38", x"E5", x"61", x"C9", x"28", x"B0", x"35",
x"C9", x"08", x"90", x"1D", x"A5", x"61", x"18", x"69",
x"08", x"85", x"61", x"A5", x"65", x"85", x"70", x"A5",
x"64", x"85", x"65", x"A5", x"63", x"85", x"64", x"A5",
x"62", x"85", x"63", x"A9", x"00", x"85", x"62", x"F0",
x"D6", x"E6", x"61", x"18", x"66", x"62", x"66", x"63",
x"66", x"64", x"66", x"65", x"66", x"70", x"A5", x"61",
x"C5", x"69", x"D0", x"ED", x"60", x"A9", x"00", x"85",
x"62", x"85", x"63", x"85", x"64", x"85", x"65", x"85",
x"70", x"A5", x"69", x"85", x"61", x"60", x"A5", x"61",
x"E5", x"69", x"C9", x"20", x"B0", x"2F", x"C9", x"08",
x"90", x"19", x"A5", x"69", x"18", x"69", x"08", x"85",
x"69", x"A5", x"6C", x"85", x"6D", x"A5", x"6B", x"85",
x"6C", x"A5", x"6A", x"85", x"6B", x"A9", x"00", x"85",
x"6A", x"F0", x"DB", x"E6", x"69", x"18", x"66", x"6A",
x"66", x"6B", x"66", x"6C", x"66", x"6D", x"A5", x"61",
x"C5", x"69", x"D0", x"EF", x"60", x"A9", x"00", x"85",
x"6A", x"85", x"6B", x"85", x"6C", x"85", x"6D", x"A5",
x"61", x"85", x"69", x"60", x"60", x"A5", x"2F", x"85",
x"47", x"A5", x"30", x"85", x"48", x"A5", x"48", x"C5",
x"32", x"D0", x"08", x"A5", x"47", x"C5", x"31", x"D0",
x"02", x"38", x"60", x"20", x"39", x"E3", x"F0", x"03",
x"4C", x"46", x"E1", x"18", x"60", x"60", x"A9", x"93",
x"20", x"D2", x"FF", x"A9", x"DA", x"A0", x"B8", x"20",
x"1E", x"AB", x"A2", x"00", x"A0", x"0A", x"20", x"0C",
x"E5", x"A9", x"C2", x"A0", x"B8", x"20", x"1E", x"AB",
x"A2", x"01", x"A0", x"0A", x"20", x"0C", x"E5", x"A2",
x"0A", x"20", x"59", x"B9", x"A9", x"55", x"A0", x"BF",
x"20", x"1E", x"AB", x"A2", x"03", x"A0", x"0A", x"20",
x"0C", x"E5", x"20", x"1E", x"A3", x"A2", x"06", x"A0",
x"00", x"20", x"0C", x"E5", x"4C", x"6B", x"A5", x"60",
x"20", x"AE", x"AD", x"A5", x"0D", x"30", x"03", x"4C",
x"C4", x"A6", x"A5", x"61", x"C9", x"06", x"F0", x"03",
x"4C", x"CC", x"A6", x"A0", x"00", x"84", x"22", x"84",
x"23", x"84", x"24", x"B1", x"62", x"20", x"F7", x"BC",
x"90", x"03", x"4C", x"CC", x"A6", x"AA", x"E0", x"00",
x"F0", x"19", x"18", x"B9", x"65", x"E2", x"65", x"22",
x"85", x"22", x"B9", x"09", x"BB", x"65", x"23", x"85",
x"23", x"B9", x"CD", x"E4", x"65", x"24", x"85", x"24",
x"CA", x"10", x"E3", x"C8", x"C0", x"06", x"D0", x"D3",
x"A4", x"24", x"A6", x"23", x"A5", x"22", x"4C", x"DB",
x"FF", x"A0", x"BF", x"A9", x"11", x"4C", x"67", x"B8",
x"20", x"25", x"E4", x"A5", x"66", x"49", x"FF", x"85",
x"66", x"4C", x"6A", x"B8", x"91", x"98", x"BF", x"B3",
x"B3", x"B1", x"4C", x"F7", x"B6", x"00", x"00", x"20",
x"25", x"E4", x"A5", x"69", x"F0", x"41", x"A5", x"61",
x"D0", x"03", x"4C", x"AD", x"A2", x"20", x"F7", x"B6",
x"A5", x"66", x"45", x"6E", x"10", x"03", x"4C", x"19",
x"A8", x"18", x"A5", x"6D", x"65", x"65", x"85", x"65",
x"A5", x"6C", x"65", x"64", x"85", x"64", x"A5", x"6B",
x"65", x"63", x"85", x"63", x"A5", x"6A", x"65", x"62",
x"85", x"62", x"B0", x"03", x"4C", x"1E", x"B5", x"E6",
x"61", x"D0", x"0D", x"A9", x"FF", x"85", x"61", x"85",
x"65", x"85", x"64", x"85", x"63", x"85", x"62", x"60",
x"38", x"66", x"62", x"66", x"63", x"66", x"64", x"66",
x"65", x"66", x"70", x"60", x"4C", x"B2", x"A6", x"4C",
x"B2", x"A6", x"4F", x"50", x"45", x"4E", x"20", x"52",
x"4F", x"4D", x"53", x"20", x"47", x"45", x"4E", x"45",
x"52", x"49", x"43", x"20", x"42", x"55", x"49", x"4C",
x"44", x"00", x"1C", x"12", x"A4", x"A4", x"A4", x"A4",
x"A4", x"A4", x"A4", x"0D", x"9E", x"12", x"A4", x"A4",
x"A4", x"A4", x"A4", x"A4", x"0D", x"1E", x"12", x"A4",
x"A4", x"A4", x"A4", x"A4", x"0D", x"9F", x"12", x"A4",
x"A4", x"A4", x"A4", x"92", x"05", x"00", x"4C", x"1E",
x"B5", x"8A", x"48", x"A5", x"62", x"85", x"25", x"A5",
x"64", x"20", x"CD", x"BC", x"85", x"22", x"86", x"23",
x"A5", x"62", x"85", x"25", x"A5", x"65", x"20", x"38",
x"B9", x"A5", x"63", x"85", x"25", x"A5", x"64", x"20",
x"38", x"B9", x"A5", x"63", x"F0", x"07", x"A5", x"65",
x"F0", x"03", x"4C", x"CA", x"A6", x"A5", x"22", x"85",
x"62", x"A5", x"23", x"85", x"63", x"68", x"AA", x"60",
x"20", x"CD", x"BC", x"E0", x"00", x"D0", x"EB", x"18",
x"65", x"23", x"B0", x"E6", x"85", x"23", x"60", x"60",
x"A5", x"52", x"C5", x"34", x"D0", x"04", x"A5", x"51",
x"C5", x"33", x"60", x"A9", x"2D", x"A0", x"B2", x"D0",
x"10", x"A9", x"D3", x"A0", x"B1", x"D0", x"0A", x"A9",
x"C0", x"A0", x"E3", x"D0", x"04", x"A9", x"8B", x"A0",
x"B0", x"20", x"DA", x"BB", x"A0", x"00", x"B1", x"35",
x"29", x"0F", x"F0", x"47", x"C9", x"0F", x"F0", x"29",
x"AA", x"BD", x"B0", x"B1", x"20", x"D2", x"FF", x"B1",
x"35", x"29", x"F0", x"F0", x"36", x"C9", x"F0", x"F0",
x"0B", x"4A", x"4A", x"4A", x"4A", x"AA", x"BD", x"B0",
x"B1", x"4C", x"9B", x"B9", x"C8", x"B1", x"35", x"AA",
x"BD", x"57", x"A2", x"20", x"D2", x"FF", x"C8", x"D0",
x"CD", x"B1", x"35", x"29", x"F0", x"BA", x"48", x"C8",
x"B1", x"35", x"29", x"0F", x"18", x"7D", x"00", x"01",
x"9A", x"AA", x"BD", x"57", x"A2", x"20", x"D2", x"FF",
x"4C", x"7F", x"B9", x"60", x"81", x"00", x"00", x"00",
x"00", x"20", x"7F", x"AF", x"C9", x"00", x"F0", x"09",
x"C9", x"3A", x"F0", x"05", x"20", x"9C", x"A6", x"18",
x"60", x"20", x"9C", x"A6", x"38", x"60", x"80", x"35",
x"04", x"F3", x"34", x"81", x"35", x"04", x"F3", x"34",
x"80", x"80", x"00", x"00", x"00", x"80", x"31", x"72",
x"17", x"F8", x"60", x"A0", x"00", x"98", x"91", x"2B",
x"C8", x"91", x"2B", x"18", x"A5", x"2B", x"69", x"02",
x"85", x"2D", x"A5", x"2C", x"69", x"00", x"85", x"2E",
x"20", x"E7", x"FF", x"A5", x"37", x"85", x"33", x"A5",
x"38", x"85", x"34", x"A5", x"2D", x"85", x"2F", x"85",
x"31", x"A5", x"2E", x"85", x"30", x"85", x"32", x"20",
x"80", x"E0", x"38", x"A5", x"2B", x"E9", x"01", x"85",
x"41", x"A5", x"2C", x"E9", x"00", x"85", x"42", x"60",
x"20", x"25", x"E4", x"4C", x"CA", x"A9", x"48", x"20",
x"7F", x"AF", x"20", x"F7", x"BC", x"B0", x"46", x"85",
x"14", x"A9", x"00", x"85", x"15", x"20", x"4D", x"A1",
x"20", x"F7", x"BC", x"B0", x"34", x"48", x"20", x"7F",
x"BA", x"B0", x"3B", x"A5", x"15", x"48", x"A5", x"14",
x"48", x"20", x"7F", x"BA", x"B0", x"2E", x"20", x"7F",
x"BA", x"B0", x"29", x"18", x"68", x"65", x"14", x"85",
x"14", x"68", x"65", x"15", x"85", x"15", x"B0", x"1E",
x"68", x"18", x"65", x"14", x"85", x"14", x"A5", x"15",
x"69", x"00", x"85", x"15", x"B0", x"11", x"4C", x"3D",
x"BA", x"20", x"9C", x"A6", x"18", x"68", x"60", x"06",
x"14", x"26", x"15", x"60", x"68", x"68", x"68", x"68",
x"AA", x"4C", x"EE", x"A6", x"4C", x"25", x"E4", x"60",
x"60", x"85", x"0A", x"20", x"59", x"F8", x"A0", x"00",
x"4C", x"BA", x"FF", x"A9", x"01", x"2C", x"A9", x"00",
x"20", x"91", x"BA", x"20", x"B5", x"E2", x"20", x"29",
x"A7", x"B0", x"08", x"20", x"8C", x"E3", x"B0", x"03",
x"20", x"9B", x"AF", x"A4", x"2C", x"A6", x"2B", x"A5",
x"0A", x"20", x"D5", x"FF", x"90", x"03", x"4C", x"AA",
x"A6", x"86", x"2D", x"84", x"2E", x"A5", x"0A", x"F0",
x"03", x"4C", x"DA", x"A1", x"20", x"00", x"BA", x"20",
x"33", x"A5", x"20", x"12", x"BC", x"A6", x"3A", x"E8",
x"D0", x"03", x"4C", x"32", x"AC", x"48", x"48", x"4C",
x"05", x"A5", x"A5", x"61", x"F0", x"0F", x"20", x"8B",
x"A4", x"20", x"87", x"AE", x"20", x"8B", x"A4", x"20",
x"8B", x"A4", x"4C", x"6A", x"B8", x"60", x"4C", x"B2",
x"A6", x"84", x"20", x"00", x"00", x"00", x"A9", x"00",
x"85", x"66", x"A0", x"BA", x"A9", x"F9", x"4C", x"0F",
x"BB", x"F5", x"4B", x"8C", x"0E", x"02", x"00", x"20",
x"25", x"E4", x"A5", x"61", x"D0", x"03", x"4C", x"C6",
x"A6", x"A5", x"69", x"D0", x"03", x"4C", x"C5", x"A9",
x"A5", x"66", x"45", x"6E", x"85", x"66", x"A9", x"A0",
x"85", x"26", x"A9", x"00", x"85", x"27", x"A5", x"69",
x"20", x"A2", x"A1", x"A5", x"26", x"38", x"E5", x"61",
x"85", x"26", x"B0", x"02", x"C6", x"27", x"A5", x"27",
x"10", x"03", x"4C", x"C5", x"A9", x"A5", x"26", x"85",
x"61", x"20", x"16", x"BF", x"20", x"95", x"A1", x"20",
x"42", x"AB", x"A5", x"6D", x"85", x"65", x"A5", x"6C",
x"85", x"64", x"A5", x"6B", x"85", x"63", x"A5", x"6A",
x"85", x"62", x"4C", x"1E", x"B5", x"A2", x"00", x"A0",
x"00", x"B1", x"35", x"C9", x"FF", x"D0", x"0A", x"C8",
x"B1", x"35", x"88", x"C9", x"FF", x"D0", x"02", x"38",
x"60", x"B1", x"35", x"D9", x"06", x"01", x"D0", x"07",
x"C9", x"00", x"F0", x"1C", x"C8", x"D0", x"F2", x"E8",
x"C9", x"00", x"F0", x"05", x"C8", x"B1", x"35", x"D0",
x"FB", x"C8", x"98", x"18", x"65", x"35", x"85", x"35",
x"A5", x"36", x"69", x"00", x"85", x"36", x"90", x"C7",
x"18", x"60", x"4C", x"9C", x"BC", x"60", x"60", x"20",
x"AE", x"AD", x"A5", x"61", x"D0", x"03", x"4C", x"BA",
x"E3", x"20", x"7F", x"AF", x"C9", x"89", x"D0", x"03",
x"4C", x"A6", x"B4", x"C9", x"A7", x"F0", x"03", x"4C",
x"CF", x"A6", x"68", x"68", x"4C", x"93", x"A4", x"4C",
x"3D", x"BC", x"4C", x"84", x"A4", x"4C", x"B2", x"A6",
x"A0", x"4A", x"A2", x"49", x"20", x"CA", x"A2", x"4C",
x"D7", x"A3", x"85", x"35", x"84", x"36", x"E0", x"00",
x"F0", x"19", x"CA", x"A0", x"00", x"B1", x"35", x"C8",
x"C9", x"00", x"D0", x"F9", x"18", x"98", x"65", x"35",
x"85", x"35", x"A9", x"00", x"65", x"36", x"85", x"36",
x"4C", x"DE", x"BB", x"60", x"4C", x"AD", x"A2", x"A5",
x"62", x"D9", x"BD", x"AA", x"D0", x"05", x"A5", x"61",
x"D9", x"A1", x"AD", x"60", x"20", x"CA", x"A2", x"4C",
x"87", x"AE", x"A5", x"2B", x"85", x"3D", x"A5", x"2C",
x"85", x"3E", x"60", x"4C", x"CA", x"A2", x"8A", x"48",
x"BA", x"E0", x"60", x"B0", x"03", x"4C", x"C1", x"A6",
x"68", x"AA", x"60", x"A5", x"61", x"F0", x"06", x"A5",
x"66", x"D0", x"02", x"A9", x"01", x"60", x"4C", x"B2",
x"A6", x"60", x"00", x"00", x"60", x"A0", x"00", x"A2",
x"57", x"4C", x"D4", x"BB", x"60", x"A9", x"00", x"85",
x"7A", x"A9", x"02", x"85", x"7B", x"A9", x"00", x"85",
x"3D", x"85", x"3E", x"A9", x"FF", x"85", x"3A", x"60",
x"60", x"00", x"00", x"60", x"A5", x"62", x"85", x"51",
x"A5", x"63", x"4C", x"6B", x"BC", x"A5", x"6A", x"85",
x"51", x"A5", x"6B", x"85", x"52", x"A2", x"19", x"E4",
x"16", x"D0", x"01", x"60", x"B4", x"00", x"F0", x"1E",
x"E8", x"B5", x"00", x"C5", x"51", x"D0", x"18", x"E8",
x"B5", x"00", x"C5", x"52", x"D0", x"12", x"84", x"50",
x"8A", x"48", x"20", x"BA", x"B3", x"68", x"AA", x"CA",
x"CA", x"A9", x"00", x"95", x"00", x"60", x"E8", x"E8",
x"E8", x"D0", x"D4", x"60", x"84", x"23", x"85", x"22",
x"A0", x"04", x"B1", x"22", x"85", x"65", x"88", x"B1",
x"22", x"85", x"64", x"88", x"B1", x"22", x"85", x"63",
x"88", x"B1", x"22", x"09", x"80", x"85", x"62", x"B1",
x"22", x"10", x"03", x"A9", x"FF", x"2C", x"A9", x"00",
x"85", x"66", x"88", x"B1", x"22", x"85", x"61", x"84",
x"70", x"A5", x"61", x"60", x"60", x"F0", x"1F", x"85",
x"24", x"A5", x"25", x"F0", x"19", x"A9", x"00", x"A2",
x"08", x"18", x"90", x"03", x"18", x"65", x"25", x"6A",
x"66", x"24", x"CA", x"10", x"F5", x"A6", x"24", x"86",
x"24", x"AA", x"A5", x"24", x"18", x"60", x"A9", x"00",
x"AA", x"18", x"60", x"60", x"4C", x"B2", x"A6", x"38",
x"E9", x"30", x"90", x"03", x"C9", x"0A", x"60", x"38",
x"60", x"20", x"95", x"B7", x"90", x"03", x"4C", x"B2",
x"A6", x"A5", x"53", x"48", x"A2", x"00", x"E8", x"20",
x"74", x"A2", x"A5", x"15", x"48", x"A5", x"14", x"48",
x"C0", x"00", x"F0", x"F2", x"86", x"61", x"20", x"23",
x"E0", x"D0", x"58", x"A9", x"05", x"20", x"D3", x"BD",
x"A9", x"00", x"85", x"62", x"85", x"63", x"A2", x"00",
x"8A", x"E8", x"0A", x"A8", x"20", x"AB", x"E0", x"20",
x"01", x"B9", x"18", x"68", x"85", x"22", x"65", x"62",
x"85", x"62", x"68", x"85", x"23", x"65", x"63", x"85",
x"63", x"A5", x"23", x"C5", x"65", x"90", x"08", x"D0",
x"2A", x"A5", x"22", x"C5", x"64", x"B0", x"24", x"E4",
x"61", x"D0", x"D5", x"68", x"85", x"53", x"85", x"64",
x"A9", x"00", x"85", x"65", x"20", x"01", x"B9", x"A5",
x"61", x"0A", x"20", x"D3", x"BD", x"18", x"A5", x"62",
x"65", x"47", x"85", x"47", x"A5", x"63", x"65", x"48",
x"85", x"48", x"60", x"4C", x"C8", x"A6", x"60", x"A9",
x"DD", x"DE", x"DF", x"E0", x"E1", x"B7", x"E2", x"F2",
x"A5", x"95", x"A6", x"19", x"E3", x"E4", x"B9", x"8F",
x"E5", x"59", x"9D", x"BD", x"9A", x"E6", x"FF", x"E7",
x"7E", x"E8", x"CB", x"FF", x"E9", x"BA", x"EA", x"EB",
x"EC", x"ED", x"ED", x"CE", x"CE", x"EE", x"A2", x"BD",
x"BD", x"BD", x"BD", x"BD", x"AE", x"BD", x"BD", x"B4",
x"B4", x"BB", x"BA", x"BD", x"BD", x"E3", x"A2", x"BD",
x"A6", x"BA", x"E2", x"BA", x"BD", x"DF", x"BD", x"BF",
x"BD", x"E3", x"B9", x"BD", x"B5", x"BD", x"BD", x"BD",
x"BF", x"BD", x"A6", x"A6", x"BD", x"4C", x"51", x"B4",
x"4C", x"B2", x"A6", x"18", x"65", x"47", x"85", x"47",
x"90", x"02", x"E6", x"48", x"60", x"60", x"EA", x"EA",
x"EA", x"EA", x"EA", x"EA", x"EA", x"EA", x"EA", x"EA",
x"EA", x"EA", x"EA", x"EA", x"EA", x"EA", x"EA", x"EA",
x"4C", x"B2", x"A6", x"20", x"46", x"A7", x"90", x"03",
x"4C", x"CF", x"A6", x"A5", x"0C", x"10", x"23", x"A9",
x"BE", x"48", x"A9", x"6B", x"48", x"A5", x"53", x"48",
x"A2", x"00", x"E8", x"20", x"74", x"A2", x"A5", x"15",
x"48", x"A5", x"14", x"48", x"C0", x"00", x"F0", x"F2",
x"8A", x"48", x"20", x"7D", x"A5", x"A9", x"FF", x"4C",
x"3F", x"BE", x"20", x"7D", x"A5", x"20", x"AD", x"AE",
x"D0", x"03", x"4C", x"F8", x"B7", x"20", x"37", x"AB",
x"D0", x"03", x"4C", x"CF", x"A6", x"20", x"66", x"BF",
x"D0", x"03", x"4C", x"CF", x"A6", x"A5", x"0C", x"48",
x"A5", x"45", x"48", x"A5", x"46", x"48", x"20", x"AE",
x"AD", x"68", x"85", x"46", x"68", x"85", x"45", x"68",
x"85", x"0C", x"10", x"23", x"A2", x"04", x"B5", x"61",
x"95", x"69", x"CA", x"10", x"F9", x"20", x"95", x"B7",
x"90", x"03", x"4C", x"B2", x"A6", x"68", x"85", x"61",
x"AA", x"4C", x"23", x"BD", x"A2", x"04", x"B5", x"69",
x"95", x"61", x"CA", x"10", x"F9", x"30", x"03", x"20",
x"AD", x"A5", x"A9", x"00", x"18", x"24", x"45", x"10",
x"02", x"69", x"01", x"24", x"46", x"10", x"02", x"69",
x"80", x"30", x"16", x"F0", x"0A", x"A5", x"0D", x"10",
x"03", x"4C", x"C4", x"A6", x"4C", x"B2", x"A6", x"A5",
x"0D", x"10", x"03", x"4C", x"C4", x"A6", x"4C", x"B2",
x"A6", x"A5", x"0D", x"30", x"03", x"4C", x"C4", x"A6",
x"20", x"EB", x"E3", x"A5", x"61", x"D0", x"0A", x"20",
x"AF", x"B3", x"A0", x"00", x"A9", x"00", x"91", x"47",
x"60", x"A5", x"51", x"C5", x"62", x"D0", x"08", x"C8",
x"A5", x"52", x"C5", x"63", x"D0", x"01", x"60", x"A5",
x"2E", x"C5", x"63", x"90", x"27", x"D0", x"06", x"A5",
x"2D", x"C5", x"62", x"90", x"1F", x"A5", x"63", x"C5",
x"2C", x"90", x"19", x"D0", x"06", x"A5", x"62", x"C5",
x"2B", x"90", x"11", x"A0", x"00", x"A5", x"61", x"91",
x"47", x"C8", x"A5", x"62", x"91", x"47", x"C8", x"A5",
x"63", x"91", x"47", x"60", x"20", x"48", x"B9", x"90",
x"0C", x"A5", x"50", x"C5", x"61", x"D0", x"03", x"4C",
x"04", x"E4", x"20", x"AF", x"B3", x"A5", x"61", x"A0",
x"00", x"91", x"47", x"20", x"D3", x"B4", x"4C", x"04",
x"E4", x"80", x"00", x"00", x"00", x"00", x"A9", x"00",
x"85", x"70", x"A5", x"65", x"D0", x"1C", x"A5", x"61",
x"C9", x"08", x"90", x"16", x"E9", x"08", x"85", x"61",
x"A5", x"64", x"85", x"65", x"A5", x"63", x"85", x"64",
x"A5", x"62", x"85", x"63", x"A9", x"00", x"85", x"62",
x"F0", x"DC", x"A5", x"65", x"29", x"01", x"D0", x"11",
x"A5", x"61", x"F0", x"0D", x"C6", x"61", x"18", x"66",
x"62", x"66", x"63", x"66", x"64", x"66", x"65", x"90",
x"E9", x"60", x"4F", x"52", x"01", x"44", x"45", x"56",
x"2E", x"32", x"30", x"31", x"32", x"30", x"36", x"2E",
x"46", x"43", x"2E", x"31", x"00", x"00", x"A5", x"46",
x"C9", x"54", x"D0", x"04", x"A5", x"45", x"C9", x"53",
x"60", x"20", x"87", x"AE", x"60", x"4C", x"B2", x"A6",
x"20", x"9C", x"BC", x"60", x"4C", x"B2", x"A6", x"20",
x"C1", x"B9", x"B0", x"2C", x"20", x"4D", x"A1", x"C9",
x"3B", x"F0", x"28", x"20", x"9C", x"A6", x"20", x"60",
x"E0", x"20", x"AE", x"AD", x"A5", x"0D", x"10", x"06",
x"20", x"44", x"E0", x"4C", x"A1", x"BF", x"4C", x"B2",
x"A6", x"20", x"C1", x"B9", x"B0", x"0A", x"C9", x"2C",
x"F0", x"E4", x"C9", x"3B", x"F0", x"05", x"D0", x"DB",
x"20", x"D2", x"F7", x"60", x"A5", x"61", x"F0", x"06",
x"A5", x"66", x"49", x"FF", x"85", x"66", x"60", x"81",
x"38", x"AA", x"3B", x"29", x"A5", x"3D", x"85", x"26",
x"A5", x"3E", x"85", x"27", x"18", x"8A", x"65", x"26",
x"85", x"24", x"A5", x"27", x"69", x"00", x"85", x"25",
x"A5", x"2D", x"38", x"E5", x"24", x"85", x"28", x"A5",
x"2E", x"E5", x"25", x"85", x"29", x"4C", x"F4", x"BF",
x"81", x"00", x"00", x"00", x"00", x"60", x"20", x"EB",
x"B9", x"4C", x"32", x"AC", x"38", x"A9", x"00", x"E5",
x"28", x"A8", x"20", x"3D", x"A2", x"4C", x"C7", x"E1",
x"20", x"2E", x"BA", x"90", x"03", x"4C", x"CF", x"A6",
x"A5", x"14", x"48", x"A5", x"15", x"48", x"20", x"C3",
x"A1", x"90", x"03", x"4C", x"CF", x"A6", x"A8", x"68",
x"85", x"15", x"68", x"85", x"14", x"98", x"A0", x"00",
x"91", x"14", x"60", x"A9", x"26", x"85", x"01", x"A0",
x"04", x"8A", x"D1", x"47", x"4C", x"B0", x"E3", x"A9",
x"26", x"85", x"01", x"A0", x"00", x"B1", x"7A", x"85",
x"3D", x"C8", x"B1", x"7A", x"85", x"3E", x"05", x"3D",
x"4C", x"B0", x"E3", x"60", x"A9", x"26", x"85", x"01",
x"A0", x"00", x"C4", x"61", x"D0", x"03", x"4C", x"61",
x"E3", x"B1", x"62", x"20", x"D2", x"FF", x"C8", x"10",
x"F1", x"60", x"4C", x"B2", x"A6", x"4C", x"B2", x"A6",
x"A2", x"19", x"E4", x"16", x"F0", x"1A", x"B5", x"00",
x"F0", x"11", x"85", x"50", x"B5", x"01", x"85", x"51",
x"B5", x"02", x"85", x"52", x"8A", x"48", x"20", x"BA",
x"B3", x"68", x"AA", x"E8", x"E8", x"E8", x"D0", x"E2",
x"A9", x"19", x"85", x"16", x"A9", x"16", x"85", x"17",
x"60", x"85", x"50", x"18", x"A5", x"22", x"65", x"50",
x"85", x"22", x"90", x"02", x"C6", x"23", x"60", x"20",
x"2B", x"BC", x"C9", x"00", x"D0", x"03", x"4C", x"22",
x"A2", x"C9", x"80", x"B0", x"03", x"4C", x"BE", x"E0",
x"4C", x"AC", x"A1", x"A9", x"26", x"85", x"01", x"B1",
x"47", x"85", x"65", x"C8", x"B1", x"47", x"85", x"64",
x"C8", x"A9", x"27", x"85", x"01", x"60", x"06", x"8C",
x"26", x"8D", x"26", x"8E", x"26", x"8F", x"B0", x"19",
x"A5", x"8C", x"49", x"B7", x"85", x"8C", x"A5", x"8D",
x"49", x"1D", x"85", x"8D", x"A5", x"8E", x"49", x"C1",
x"85", x"8E", x"A5", x"8F", x"49", x"04", x"85", x"8F",
x"38", x"A5", x"8E", x"69", x"C6", x"85", x"62", x"A5",
x"8C", x"49", x"4E", x"85", x"63", x"A5", x"8F", x"49",
x"62", x"85", x"64", x"A5", x"8D", x"24", x"8D", x"2A",
x"85", x"65", x"A9", x"00", x"85", x"66", x"A9", x"80",
x"85", x"70", x"85", x"61", x"4C", x"1E", x"B5", x"AA",
x"A5", x"16", x"C9", x"22", x"B0", x"13", x"A8", x"85",
x"17", x"18", x"69", x"03", x"85", x"16", x"96", x"00",
x"84", x"47", x"A9", x"00", x"85", x"48", x"4C", x"D3",
x"B4", x"A0", x"19", x"B9", x"00", x"00", x"F0", x"EE",
x"C8", x"C8", x"C8", x"C0", x"22", x"D0", x"F4", x"4C",
x"C1", x"A6", x"A9", x"26", x"85", x"01", x"A0", x"00",
x"B1", x"3D", x"48", x"C8", x"B1", x"3D", x"85", x"3E",
x"68", x"85", x"3D", x"4C", x"61", x"E3", x"A9", x"26",
x"85", x"01", x"A0", x"03", x"B1", x"47", x"48", x"88",
x"B1", x"47", x"18", x"65", x"47", x"85", x"47", x"68",
x"65", x"48", x"85", x"48", x"A9", x"27", x"85", x"01",
x"4C", x"9D", x"B7", x"A9", x"26", x"85", x"01", x"A0",
x"00", x"B1", x"22", x"F0", x"18", x"C8", x"18", x"71",
x"22", x"85", x"26", x"C8", x"A9", x"00", x"71", x"22",
x"85", x"27", x"A0", x"00", x"A5", x"22", x"91", x"26",
x"C8", x"A5", x"23", x"91", x"26", x"4C", x"61", x"E3",
x"A9", x"26", x"85", x"01", x"B1", x"7A", x"48", x"A9",
x"27", x"85", x"01", x"68", x"60", x"A9", x"26", x"85",
x"01", x"B1", x"3D", x"4C", x"8E", x"E1", x"A9", x"26",
x"85", x"01", x"B1", x"47", x"4C", x"8E", x"E1", x"A9",
x"26", x"85", x"01", x"B1", x"62", x"4C", x"8E", x"E1",
x"08", x"A9", x"26", x"85", x"01", x"B1", x"24", x"91",
x"26", x"88", x"D0", x"F9", x"C6", x"25", x"C6", x"27",
x"C6", x"29", x"D0", x"F1", x"4C", x"DB", x"E1", x"08",
x"A9", x"26", x"85", x"01", x"B1", x"24", x"91", x"26",
x"C8", x"D0", x"F9", x"E6", x"25", x"E6", x"27", x"C6",
x"29", x"D0", x"F1", x"A9", x"27", x"85", x"01", x"28",
x"60", x"A9", x"26", x"85", x"01", x"A0", x"02", x"B1",
x"22", x"18", x"65", x"22", x"85", x"24", x"C8", x"B1",
x"22", x"65", x"23", x"85", x"25", x"A0", x"00", x"B1",
x"22", x"10", x"03", x"4C", x"5E", x"E2", x"C8", x"B1",
x"22", x"30", x"03", x"4C", x"5E", x"E2", x"A0", x"04",
x"B1", x"22", x"0A", x"18", x"69", x"05", x"20", x"89",
x"E0", x"4C", x"58", x"E2", x"20", x"12", x"BC", x"A9",
x"26", x"85", x"01", x"20", x"4C", x"E2", x"F0", x"3E",
x"A0", x"03", x"B1", x"3D", x"C5", x"15", x"F0", x"04",
x"B0", x"34", x"D0", x"0B", x"88", x"B1", x"3D", x"C5",
x"14", x"F0", x"25", x"B0", x"29", x"D0", x"00", x"20",
x"4C", x"E2", x"F0", x"22", x"A0", x"00", x"B1", x"3D",
x"48", x"C8", x"B1", x"3D", x"85", x"3E", x"68", x"85",
x"3D", x"4C", x"17", x"E2", x"A0", x"01", x"B1", x"3D",
x"D0", x"05", x"88", x"B1", x"3D", x"D0", x"00", x"60",
x"A9", x"27", x"85", x"01", x"18", x"60", x"A9", x"27",
x"85", x"01", x"38", x"60", x"60", x"80", x"C0", x"A0",
x"10", x"58", x"3C", x"60", x"05", x"67", x"CC", x"65",
x"20", x"E2", x"6E", x"38", x"AD", x"08", x"B4", x"74",
x"D0", x"0B", x"7B", x"30", x"7A", x"08", x"88", x"84",
x"2A", x"7E", x"AA", x"AA", x"AA", x"95", x"81", x"00",
x"00", x"00", x"00", x"CE", x"01", x"01", x"CE", x"01",
x"01", x"38", x"A5", x"07", x"ED", x"01", x"01", x"85",
x"07", x"EE", x"00", x"01", x"AC", x"00", x"01", x"AD",
x"01", x"01", x"18", x"6D", x"00", x"01", x"AA", x"BD",
x"00", x"02", x"99", x"00", x"02", x"F0", x"04", x"E8",
x"C8", x"D0", x"F4", x"60", x"60", x"A9", x"01", x"A2",
x"41", x"A0", x"F1", x"4C", x"BD", x"FF", x"20", x"93",
x"BA", x"20", x"29", x"A7", x"90", x"03", x"4C", x"D2",
x"A6", x"20", x"8C", x"E3", x"B0", x"03", x"20", x"9B",
x"AF", x"A9", x"2B", x"A6", x"2D", x"A4", x"2E", x"20",
x"D8", x"FF", x"90", x"03", x"4C", x"AA", x"A6", x"60",
x"81", x"49", x"0F", x"DA", x"A2", x"83", x"49", x"0F",
x"DA", x"A2", x"7F", x"00", x"00", x"00", x"00", x"EA",
x"EA", x"EA", x"EA", x"EA", x"EA", x"EA", x"EA", x"EA",
x"EA", x"EA", x"EA", x"EA", x"EA", x"EA", x"EA", x"EA",
x"EA", x"EA", x"EA", x"EA", x"EA", x"EA", x"4C", x"B2",
x"A6", x"83", x"49", x"0F", x"DA", x"A2", x"60", x"4C",
x"B2", x"A6", x"A5", x"2B", x"85", x"3D", x"A5", x"2C",
x"85", x"3E", x"A5", x"3D", x"85", x"2D", x"A5", x"3E",
x"85", x"2E", x"20", x"32", x"E1", x"A5", x"3D", x"05",
x"3E", x"D0", x"EF", x"18", x"A5", x"2D", x"69", x"02",
x"85", x"2D", x"90", x"02", x"E6", x"2E", x"4C", x"00",
x"BA", x"A9", x"26", x"85", x"01", x"A0", x"00", x"B1",
x"47", x"C5", x"45", x"D0", x"05", x"C8", x"B1", x"47",
x"C5", x"46", x"4C", x"B0", x"E3", x"A9", x"26", x"85",
x"01", x"A0", x"00", x"B1", x"47", x"85", x"61", x"C8",
x"B1", x"47", x"85", x"62", x"C8", x"B1", x"47", x"85",
x"63", x"A9", x"27", x"85", x"01", x"60", x"A9", x"26",
x"85", x"01", x"B1", x"3D", x"85", x"24", x"C8", x"B1",
x"3D", x"85", x"25", x"4C", x"88", x"E3", x"A9", x"26",
x"85", x"01", x"B1", x"3D", x"18", x"65", x"22", x"91",
x"3D", x"C8", x"B1", x"3D", x"65", x"23", x"91", x"3D",
x"4C", x"61", x"E3", x"60", x"20", x"C3", x"A1", x"B0",
x"02", x"85", x"BA", x"60", x"A0", x"13", x"B9", x"52",
x"BF", x"D9", x"B9", x"E4", x"F0", x"05", x"A9", x"01",
x"6C", x"B7", x"E4", x"88", x"10", x"F0", x"4C", x"E5",
x"A7", x"A9", x"26", x"85", x"01", x"20", x"4C", x"E2",
x"08", x"A9", x"27", x"85", x"01", x"28", x"60", x"4C",
x"F1", x"A1", x"48", x"48", x"4C", x"E9", x"A4", x"60",
x"4B", x"FA", x"0F", x"00", x"83", x"EB", x"00", x"4A",
x"05", x"00", x"FF", x"FF", x"20", x"12", x"BC", x"A0",
x"01", x"20", x"95", x"E1", x"C9", x"00", x"D0", x"03",
x"4C", x"32", x"AC", x"A5", x"91", x"30", x"03", x"4C",
x"90", x"A2", x"20", x"85", x"AB", x"20", x"32", x"E1",
x"4C", x"CF", x"E3", x"A9", x"26", x"85", x"01", x"A0",
x"00", x"B1", x"47", x"85", x"50", x"C8", x"B1", x"47",
x"85", x"51", x"C8", x"B1", x"47", x"85", x"52", x"A9",
x"27", x"85", x"01", x"60", x"A9", x"26", x"85", x"01",
x"A0", x"02", x"B1", x"47", x"85", x"52", x"88", x"B1",
x"47", x"85", x"51", x"88", x"B1", x"62", x"91", x"51",
x"C8", x"C4", x"61", x"D0", x"F7", x"A9", x"27", x"85",
x"01", x"60", x"4C", x"B6", x"B7", x"84", x"23", x"85",
x"22", x"A0", x"04", x"B1", x"22", x"85", x"6D", x"88",
x"B1", x"22", x"85", x"6C", x"88", x"B1", x"22", x"85",
x"6B", x"88", x"B1", x"22", x"09", x"80", x"85", x"6A",
x"B1", x"22", x"10", x"03", x"A9", x"FF", x"2C", x"A9",
x"00", x"85", x"6E", x"88", x"B1", x"22", x"85", x"69",
x"A5", x"61", x"60", x"60", x"4C", x"B2", x"A6", x"38",
x"A5", x"2D", x"E9", x"01", x"85", x"24", x"A5", x"2E",
x"E9", x"00", x"85", x"25", x"18", x"8A", x"65", x"24",
x"85", x"26", x"A5", x"25", x"69", x"00", x"85", x"27",
x"A5", x"2D", x"38", x"E5", x"3D", x"85", x"28", x"A5",
x"2E", x"E5", x"3E", x"85", x"29", x"4C", x"A6", x"AD",
x"A9", x"26", x"85", x"01", x"B1", x"3D", x"85", x"39",
x"C8", x"B1", x"3D", x"85", x"3A", x"A9", x"27", x"85",
x"01", x"4C", x"93", x"A4", x"A9", x"26", x"85", x"01",
x"A0", x"00", x"B1", x"6A", x"91", x"22", x"C8", x"C4",
x"69", x"D0", x"F7", x"98", x"20", x"89", x"E0", x"A0",
x"00", x"B1", x"62", x"91", x"22", x"C8", x"C4", x"61",
x"D0", x"F7", x"A9", x"27", x"85", x"01", x"60", x"54",
x"ED", x"4F", x"52", x"01", x"44", x"45", x"56", x"2E",
x"32", x"30", x"31", x"32", x"30", x"36", x"2E", x"46",
x"43", x"2E", x"31", x"00", x"00", x"20", x"03", x"00",
x"00", x"00", x"00", x"E6", x"A2", x"D0", x"06", x"E6",
x"A1", x"D0", x"02", x"E6", x"A0", x"A5", x"A0", x"C9",
x"4F", x"90", x"0E", x"A5", x"A1", x"C9", x"1A", x"90",
x"08", x"A9", x"00", x"85", x"A0", x"85", x"A1", x"85",
x"A2", x"A9", x"80", x"8D", x"00", x"DC", x"AD", x"01",
x"DC", x"49", x"FF", x"85", x"91", x"A9", x"7F", x"8D",
x"00", x"DC", x"AD", x"01", x"DC", x"05", x"91", x"85",
x"91", x"60", x"B0", x"07", x"84", x"D3", x"86", x"D6",
x"20", x"6C", x"E5", x"A4", x"D3", x"A6", x"D6", x"60",
x"20", x"A0", x"E5", x"4C", x"20", x"FC", x"85", x"9D",
x"60", x"B9", x"59", x"02", x"D0", x"03", x"4C", x"7B",
x"F2", x"B9", x"63", x"02", x"20", x"6A", x"F9", x"90",
x"03", x"4C", x"87", x"EA", x"B9", x"59", x"02", x"09",
x"60", x"20", x"B7", x"E6", x"90", x"03", x"4C", x"87",
x"EA", x"4C", x"73", x"F2", x"A9", x"80", x"A0", x"18",
x"99", x"D9", x"00", x"88", x"10", x"FA", x"A2", x"18",
x"20", x"FF", x"E9", x"CA", x"10", x"FA", x"4C", x"66",
x"E5", x"20", x"94", x"E5", x"90", x"03", x"4C", x"79",
x"FC", x"09", x"E0", x"4C", x"89", x"E5", x"A9", x"00",
x"85", x"D3", x"85", x"D6", x"20", x"E6", x"EB", x"4C",
x"B6", x"FC", x"20", x"94", x"E5", x"90", x"03", x"4C",
x"79", x"FC", x"09", x"F0", x"85", x"A4", x"20", x"DA",
x"FA", x"B0", x"10", x"20", x"61", x"FF", x"4C", x"CD",
x"F4", x"85", x"A4", x"20", x"DA", x"FA", x"B0", x"03",
x"4C", x"CD", x"F4", x"60", x"C9", x"10", x"90", x"06",
x"C9", x"60", x"F0", x"02", x"38", x"60", x"18", x"60",
x"A9", x"00", x"A2", x"2E", x"9D", x"00", x"D0", x"CA",
x"10", x"FA", x"A9", x"1B", x"8D", x"11", x"D0", x"A9",
x"C8", x"8D", x"16", x"D0", x"A9", x"14", x"8D", x"18",
x"D0", x"A9", x"0F", x"8D", x"19", x"D0", x"A9", x"06",
x"8D", x"20", x"D0", x"8D", x"21", x"D0", x"4C", x"36",
x"F3", x"A0", x"19", x"A2", x"28", x"60", x"68", x"68",
x"58", x"4C", x"67", x"FC", x"A5", x"01", x"29", x"10",
x"F0", x"10", x"A2", x"35", x"20", x"50", x"F9", x"20",
x"ED", x"F6", x"B0", x"EA", x"A5", x"01", x"29", x"10",
x"D0", x"F5", x"A9", x"01", x"85", x"C0", x"A2", x"4F",
x"20", x"50", x"F9", x"20", x"D2", x"F7", x"4C", x"9D",
x"FB", x"20", x"92", x"FB", x"A2", x"49", x"20", x"50",
x"F9", x"A0", x"05", x"B1", x"B2", x"20", x"D2", x"FF",
x"C8", x"C0", x"15", x"D0", x"F6", x"20", x"8A", x"E6",
x"B0", x"BC", x"20", x"65", x"E6", x"B0", x"46", x"A0",
x"01", x"B1", x"B2", x"85", x"C1", x"C8", x"B1", x"B2",
x"85", x"C2", x"C8", x"B1", x"B2", x"85", x"AE", x"C8",
x"B1", x"B2", x"85", x"AF", x"A5", x"B9", x"D0", x"22",
x"38", x"A5", x"AE", x"E5", x"C1", x"85", x"AE", x"A5",
x"AF", x"E5", x"C2", x"85", x"AF", x"A5", x"C3", x"85",
x"C1", x"A5", x"C4", x"85", x"C2", x"18", x"A5", x"AE",
x"65", x"C1", x"85", x"AE", x"A5", x"AF", x"65", x"C2",
x"85", x"AF", x"20", x"B0", x"FE", x"20", x"E5", x"FE",
x"20", x"9D", x"FB", x"18", x"60", x"20", x"D2", x"F7",
x"20", x"9D", x"FB", x"38", x"60", x"A5", x"B7", x"F0",
x"F2", x"A0", x"00", x"A9", x"20", x"C4", x"B7", x"B0",
x"02", x"B1", x"BB", x"C9", x"2A", x"F0", x"E4", x"C8",
x"C8", x"C8", x"C8", x"C8", x"D1", x"B2", x"D0", x"E3",
x"88", x"88", x"88", x"88", x"C0", x"10", x"D0", x"E3",
x"18", x"60", x"A0", x"00", x"20", x"F1", x"E4", x"A5",
x"91", x"10", x"12", x"29", x"10", x"F0", x"0C", x"A2",
x"80", x"20", x"8D", x"F9", x"CA", x"20", x"8D", x"F9",
x"88", x"D0", x"E9", x"18", x"60", x"38", x"60", x"20",
x"92", x"FB", x"20", x"17", x"FF", x"4C", x"3D", x"FF",
x"20", x"92", x"FB", x"4C", x"4F", x"FF", x"60", x"4C",
x"89", x"E5", x"78", x"A0", x"00", x"AD", x"00", x"DD",
x"29", x"C7", x"85", x"A3", x"09", x"20", x"85", x"A4",
x"2C", x"00", x"DD", x"50", x"FB", x"A5", x"A3", x"8D",
x"00", x"DD", x"A2", x"13", x"2C", x"00", x"DD", x"50",
x"16", x"CA", x"D0", x"F8", x"20", x"9D", x"FA", x"AD",
x"01", x"DD", x"91", x"AE", x"38", x"20", x"76", x"F8",
x"A9", x"02", x"85", x"A3", x"4C", x"DF", x"E7", x"AD",
x"01", x"DD", x"91", x"AE", x"A5", x"A4", x"8D", x"00",
x"DD", x"C8", x"D0", x"CC", x"E6", x"AF", x"4C", x"C8",
x"E6", x"60", x"AD", x"12", x"D0", x"C9", x"2E", x"90",
x"0C", x"AD", x"12", x"D0", x"ED", x"11", x"D0", x"29",
x"07", x"C9", x"06", x"B0", x"F4", x"60", x"60", x"AD",
x"00", x"DD", x"29", x"07", x"85", x"94", x"60", x"C9",
x"E0", x"B0", x"07", x"C9", x"C0", x"90", x"03", x"29",
x"7F", x"60", x"C9", x"40", x"90", x"0E", x"38", x"E9",
x"40", x"C9", x"20", x"90", x"07", x"C9", x"40", x"B0",
x"03", x"18", x"69", x"20", x"60", x"4C", x"43", x"FF",
x"4C", x"73", x"FC", x"A5", x"BA", x"20", x"24", x"FA",
x"4C", x"4F", x"FF", x"68", x"A5", x"BA", x"20", x"24",
x"FA", x"4C", x"67", x"FC", x"A5", x"B7", x"D0", x"03",
x"4C", x"7F", x"FC", x"20", x"CB", x"FE", x"A5", x"BA",
x"20", x"6A", x"F9", x"B0", x"D8", x"A9", x"00", x"20",
x"72", x"E5", x"B0", x"D1", x"20", x"5C", x"FB", x"B0",
x"D2", x"A5", x"BA", x"20", x"66", x"FA", x"B0", x"CB",
x"A9", x"60", x"85", x"A4", x"20", x"DA", x"FA", x"B0",
x"C2", x"20", x"61", x"FF", x"20", x"AD", x"FB", x"B0",
x"BA", x"20", x"EA", x"E7", x"85", x"AE", x"20", x"EA",
x"E7", x"85", x"AF", x"A5", x"B9", x"D0", x"08", x"A5",
x"C1", x"85", x"AE", x"A5", x"C2", x"85", x"AF", x"20",
x"E5", x"FE", x"A5", x"93", x"D0", x"10", x"A5", x"A3",
x"C9", x"01", x"D0", x"03", x"4C", x"7D", x"EF", x"C9",
x"02", x"D0", x"03", x"4C", x"BA", x"E6", x"20", x"21",
x"EF", x"B0", x"88", x"20", x"99", x"FE", x"B0", x"83",
x"E6", x"AE", x"D0", x"02", x"E6", x"AF", x"A5", x"AE",
x"29", x"1F", x"D0", x"0F", x"8A", x"48", x"20", x"F1",
x"E4", x"20", x"ED", x"F6", x"90", x"03", x"4C", x"4B",
x"E7", x"68", x"AA", x"24", x"90", x"50", x"D7", x"20",
x"17", x"FF", x"A5", x"BA", x"20", x"24", x"FA", x"4C",
x"3D", x"FF", x"20", x"21", x"EF", x"B0", x"09", x"A5",
x"90", x"29", x"40", x"D0", x"03", x"A5", x"A4", x"60",
x"68", x"68", x"4C", x"40", x"E7", x"AD", x"8D", x"02",
x"8D", x"8E", x"02", x"A9", x"00", x"8D", x"8D", x"02",
x"A2", x"00", x"8E", x"00", x"DC", x"CA", x"EC", x"01",
x"DC", x"F0", x"72", x"A0", x"03", x"B9", x"D7", x"F8",
x"8D", x"00", x"DC", x"B9", x"DB", x"F8", x"2D", x"01",
x"DC", x"D0", x"09", x"AD", x"8D", x"02", x"19", x"DF",
x"F8", x"8D", x"8D", x"02", x"88", x"10", x"E6", x"AD",
x"90", x"02", x"D0", x"06", x"20", x"48", x"EB", x"4C",
x"3D", x"E8", x"20", x"69", x"F1", x"20", x"DC", x"F7",
x"EC", x"01", x"DC", x"D0", x"40", x"A5", x"F6", x"F0",
x"3C", x"A0", x"FF", x"A2", x"07", x"BD", x"16", x"F8",
x"8D", x"00", x"DC", x"BD", x"36", x"F8", x"0D", x"01",
x"DC", x"C9", x"FF", x"F0", x"19", x"C0", x"FF", x"D0",
x"24", x"A0", x"07", x"D9", x"16", x"F8", x"D0", x"09",
x"98", x"18", x"7D", x"26", x"F8", x"A8", x"4C", x"76",
x"E8", x"88", x"10", x"EF", x"30", x"0F", x"CA", x"10",
x"D4", x"C0", x"FF", x"F0", x"08", x"20", x"DC", x"F7",
x"EC", x"01", x"DC", x"F0", x"05", x"A9", x"40", x"85",
x"C5", x"60", x"C4", x"C5", x"F0", x"1F", x"84", x"C5",
x"A9", x"16", x"8D", x"8C", x"02", x"A5", x"C6", x"CD",
x"89", x"02", x"B0", x"35", x"A9", x"03", x"8D", x"8B",
x"02", x"B1", x"F5", x"F0", x"E0", x"A4", x"C6", x"99",
x"77", x"02", x"E6", x"C6", x"60", x"AD", x"8A", x"02",
x"30", x"0D", x"98", x"A2", x"03", x"DD", x"F7", x"F3",
x"F0", x"05", x"CA", x"10", x"F8", x"30", x"ED", x"AD",
x"8C", x"02", x"F0", x"04", x"CE", x"8C", x"02", x"60",
x"AD", x"8B", x"02", x"F0", x"C8", x"CE", x"8B", x"02",
x"60", x"A9", x"00", x"8D", x"8C", x"02", x"8D", x"8B",
x"02", x"60", x"90", x"05", x"1C", x"9F", x"9C", x"1E",
x"1F", x"9E", x"81", x"95", x"96", x"97", x"98", x"99",
x"9A", x"9B", x"AD", x"8D", x"02", x"29", x"04", x"F0",
x"0A", x"A0", x"09", x"A2", x"FF", x"20", x"8D", x"F9",
x"88", x"D0", x"F8", x"A0", x"00", x"B9", x"DA", x"00",
x"99", x"D9", x"00", x"C8", x"C0", x"18", x"D0", x"F5",
x"A9", x"80", x"85", x"F1", x"20", x"FA", x"F9", x"AD",
x"88", x"02", x"85", x"AD", x"85", x"AF", x"A9", x"D8",
x"85", x"D2", x"85", x"F4", x"A9", x"00", x"85", x"AE",
x"85", x"F3", x"A9", x"28", x"85", x"AC", x"85", x"D1",
x"A0", x"00", x"B1", x"AC", x"91", x"AE", x"B1", x"D1",
x"91", x"F3", x"C0", x"BF", x"D0", x"06", x"A5", x"F4",
x"C9", x"DB", x"F0", x"0D", x"C8", x"D0", x"EB", x"E6",
x"AD", x"E6", x"AF", x"E6", x"F4", x"E6", x"D2", x"D0",
x"E1", x"20", x"34", x"FE", x"A2", x"18", x"20", x"FF",
x"E9", x"C6", x"D6", x"24", x"D9", x"10", x"93", x"4C",
x"E6", x"EB", x"8A", x"48", x"A9", x"01", x"85", x"A7",
x"20", x"41", x"FB", x"26", x"A7", x"90", x"F9", x"68",
x"AA", x"A5", x"A7", x"60", x"60", x"2C", x"00", x"DD",
x"50", x"FB", x"60", x"86", x"97", x"98", x"48", x"A5",
x"D0", x"F0", x"25", x"C5", x"C8", x"D0", x"0E", x"A9",
x"00", x"85", x"D0", x"85", x"D4", x"68", x"A8", x"A6",
x"97", x"18", x"A9", x"0D", x"60", x"E6", x"D0", x"A8",
x"B1", x"C9", x"20", x"09", x"F9", x"AA", x"68", x"A8",
x"8A", x"A6", x"97", x"20", x"43", x"EC", x"18", x"60",
x"20", x"CD", x"F7", x"A5", x"C6", x"F0", x"D0", x"AD",
x"77", x"02", x"C9", x"0D", x"D0", x"40", x"20", x"C1",
x"ED", x"20", x"1D", x"FD", x"20", x"C5", x"ED", x"A5",
x"D1", x"85", x"C9", x"A5", x"D2", x"85", x"CA", x"A4",
x"D6", x"B9", x"D9", x"00", x"30", x"0F", x"A5", x"C9",
x"38", x"E9", x"28", x"85", x"C9", x"B0", x"02", x"C6",
x"CA", x"A0", x"50", x"D0", x"04", x"20", x"50", x"FA",
x"C8", x"88", x"30", x"A9", x"B1", x"C9", x"C9", x"20",
x"F0", x"F7", x"C8", x"84", x"C8", x"A0", x"01", x"84",
x"D0", x"88", x"84", x"D4", x"F0", x"A2", x"AD", x"77",
x"02", x"20", x"C9", x"FB", x"90", x"B8", x"20", x"CA",
x"F1", x"20", x"1D", x"FD", x"4C", x"77", x"E9", x"8A",
x"48", x"20", x"E8", x"EB", x"68", x"AA", x"A0", x"27",
x"AD", x"86", x"02", x"91", x"F3", x"A9", x"20", x"91",
x"D1", x"88", x"10", x"F4", x"60", x"A9", x"06", x"8D",
x"20", x"D0", x"20", x"19", x"FA", x"B0", x"10", x"20",
x"74", x"EC", x"B0", x"0B", x"C4", x"A7", x"D0", x"07",
x"88", x"29", x"7E", x"D0", x"E8", x"18", x"60", x"38",
x"60", x"20", x"9A", x"ED", x"20", x"9F", x"FF", x"20",
x"EA", x"FF", x"A5", x"01", x"29", x"10", x"F0", x"09",
x"20", x"EF", x"F8", x"A9", x"00", x"85", x"C0", x"F0",
x"07", x"A5", x"C0", x"D0", x"03", x"20", x"F5", x"F8",
x"4C", x"7E", x"EA", x"48", x"8A", x"48", x"98", x"48",
x"D8", x"BA", x"BD", x"04", x"01", x"29", x"10", x"D0",
x"0B", x"AD", x"15", x"03", x"F0", x"03", x"6C", x"14",
x"03", x"4C", x"31", x"EA", x"38", x"BD", x"05", x"01",
x"E9", x"02", x"85", x"B0", x"BD", x"06", x"01", x"E9",
x"00", x"85", x"B1", x"6C", x"16", x"03", x"AC", x"0D",
x"DC", x"68", x"A8", x"68", x"AA", x"68", x"40", x"68",
x"A8", x"68", x"20", x"A6", x"F9", x"4C", x"76", x"FC",
x"68", x"A8", x"68", x"4C", x"70", x"FC", x"A9", x"0B",
x"8D", x"20", x"D0", x"A9", x"00", x"8D", x"18", x"D4",
x"A9", x"00", x"85", x"97", x"A0", x"60", x"20", x"91",
x"FD", x"20", x"91", x"FD", x"C9", x"28", x"90", x"F0",
x"C9", x"E8", x"B0", x"EC", x"C9", x"B9", x"90", x"02",
x"C6", x"97", x"C9", x"97", x"B0", x"02", x"E6", x"97",
x"A5", x"97", x"C9", x"FD", x"F0", x"09", x"88", x"10",
x"E0", x"A5", x"97", x"30", x"02", x"18", x"60", x"38",
x"60", x"0D", x"53", x"45", x"41", x"52", x"43", x"48",
x"49", x"4E", x"47", x"20", x"46", x"4F", x"52", x"A0",
x"0D", x"4C", x"4F", x"41", x"44", x"49", x"4E", x"C7",
x"0D", x"56", x"45", x"52", x"49", x"46", x"59", x"49",
x"4E", x"C7", x"0D", x"53", x"41", x"56", x"49", x"4E",
x"47", x"A0", x"20", x"46", x"52", x"4F", x"4D", x"20",
x"A4", x"20", x"54", x"4F", x"20", x"A4", x"0D", x"50",
x"52", x"45", x"53", x"53", x"20", x"50", x"4C", x"41",
x"59", x"20", x"4F", x"4E", x"20", x"54", x"41", x"50",
x"45", x"8D", x"46", x"4F", x"55", x"4E", x"44", x"A0",
x"4F", x"4B", x"0D", x"0D", x"53", x"45", x"41", x"52",
x"43", x"48", x"49", x"4E", x"C7", x"4B", x"45", x"52",
x"4E", x"41", x"4C", x"20", x"50", x"41", x"4E", x"49",
x"C3", x"20", x"2D", x"20", x"52", x"4F", x"4D", x"20",
x"4D", x"49", x"53", x"4D", x"41", x"54", x"43", x"C8",
x"A9", x"DD", x"85", x"F5", x"A9", x"F4", x"85", x"F6",
x"AD", x"8D", x"02", x"29", x"07", x"AA", x"BD", x"2E",
x"F8", x"C9", x"FF", x"D0", x"04", x"A9", x"00", x"F0",
x"09", x"18", x"65", x"F5", x"85", x"F5", x"A9", x"00",
x"65", x"F6", x"85", x"F6", x"AD", x"91", x"02", x"D0",
x"1A", x"AD", x"8D", x"02", x"29", x"03", x"C9", x"03",
x"D0", x"11", x"AD", x"8E", x"02", x"29", x"03", x"C9",
x"03", x"F0", x"08", x"AD", x"18", x"D0", x"49", x"02",
x"8D", x"18", x"D0", x"60", x"20", x"44", x"E5", x"4C",
x"22", x"EE", x"A5", x"01", x"48", x"29", x"FE", x"85",
x"01", x"B1", x"C3", x"AA", x"68", x"85", x"01", x"8A",
x"60", x"A5", x"01", x"48", x"29", x"FE", x"85", x"01",
x"B1", x"BB", x"4C", x"9B", x"EB", x"A5", x"01", x"48",
x"29", x"FE", x"85", x"01", x"B1", x"AE", x"4C", x"9B",
x"EB", x"83", x"85", x"89", x"86", x"8A", x"87", x"88",
x"5F", x"4C", x"00", x"40", x"38", x"24", x"00", x"4C",
x"4F", x"41", x"44", x"00", x"40", x"39", x"24", x"00",
x"52", x"55", x"4E", x"3A", x"00", x"40", x"31", x"30",
x"24", x"00", x"40", x"31", x"31", x"24", x"00", x"00",
x"03", x"07", x"0C", x"10", x"15", x"1A", x"A6", x"D6",
x"AD", x"88", x"02", x"85", x"D2", x"A9", x"00", x"85",
x"D1", x"E0", x"00", x"F0", x"0E", x"A9", x"28", x"18",
x"65", x"D1", x"85", x"D1", x"90", x"02", x"E6", x"D2",
x"CA", x"D0", x"F2", x"A5", x"D1", x"85", x"F3", x"A5",
x"D2", x"38", x"ED", x"88", x"02", x"18", x"69", x"D8",
x"85", x"F4", x"60", x"93", x"13", x"08", x"09", x"0E",
x"8E", x"92", x"12", x"1D", x"9D", x"11", x"91", x"94",
x"03", x"14", x"0D", x"8B", x"F3", x"A1", x"9E", x"B7",
x"AC", x"6E", x"6B", x"BE", x"CD", x"B0", x"A7", x"FC",
x"3D", x"8C", x"76", x"EB", x"F7", x"F8", x"F8", x"F9",
x"F9", x"F8", x"F8", x"EC", x"EC", x"EC", x"EC", x"F5",
x"F8", x"F3", x"FB", x"C9", x"20", x"90", x"1F", x"C9",
x"40", x"90", x"1D", x"C9", x"60", x"90", x"1A", x"C9",
x"80", x"90", x"13", x"24", x"D4", x"30", x"15", x"C9",
x"A0", x"90", x"16", x"C9", x"C0", x"90", x"0A", x"C9",
x"E0", x"90", x"05", x"18", x"90", x"0B", x"69", x"40",
x"60", x"69", x"80", x"60", x"C9", x"C0", x"90", x"F9",
x"18", x"69", x"C0", x"60", x"A9", x"01", x"85", x"9B",
x"A9", x"7F", x"85", x"A7", x"20", x"E6", x"FB", x"B0",
x"22", x"F0", x"07", x"A9", x"01", x"45", x"9B", x"85",
x"9B", x"38", x"66", x"A7", x"B0", x"EE", x"20", x"E6",
x"FB", x"B0", x"10", x"F0", x"02", x"A9", x"01", x"45",
x"9B", x"D0", x"08", x"A2", x"0B", x"8E", x"20", x"D0",
x"A5", x"A7", x"60", x"A2", x"09", x"38", x"B0", x"F5",
x"A5", x"D6", x"F0", x"02", x"C6", x"D6", x"4C", x"22",
x"EE", x"A5", x"D6", x"C9", x"18", x"D0", x"03", x"20",
x"EA", x"E8", x"E6", x"D6", x"4C", x"22", x"EE", x"20",
x"FC", x"F8", x"C0", x"27", x"D0", x"03", x"4C", x"BF",
x"F9", x"C8", x"84", x"D3", x"10", x"E0", x"20", x"FC",
x"F8", x"88", x"10", x"F6", x"A5", x"D6", x"F0", x"D6",
x"C6", x"D6", x"A9", x"27", x"85", x"D3", x"D0", x"CE",
x"A9", x"BF", x"85", x"92", x"20", x"27", x"FB", x"B0",
x"30", x"A2", x"C0", x"A0", x"04", x"86", x"97", x"20",
x"5A", x"E9", x"C9", x"02", x"D0", x"EA", x"88", x"D0",
x"F4", x"A6", x"97", x"CA", x"D0", x"ED", x"20", x"27",
x"FB", x"B0", x"16", x"A2", x"09", x"20", x"5A", x"E9",
x"C9", x"02", x"F0", x"F9", x"A0", x"00", x"E4", x"A7",
x"D0", x"EC", x"20", x"5A", x"E9", x"CA", x"D0", x"F6",
x"18", x"60", x"A9", x"91", x"85", x"92", x"A9", x"67",
x"85", x"96", x"A9", x"80", x"A0", x"FF", x"30", x"07",
x"A9", x"04", x"2C", x"A9", x"01", x"A0", x"00", x"84",
x"A7", x"85", x"BE", x"A9", x"0B", x"8D", x"20", x"D0",
x"A5", x"BE", x"85", x"BD", x"A0", x"40", x"20", x"91",
x"FD", x"90", x"F5", x"24", x"A7", x"10", x"04", x"C9",
x"B9", x"B0", x"08", x"88", x"D0", x"F0", x"C6", x"BD",
x"D0", x"EA", x"18", x"60", x"48", x"78", x"20", x"A3",
x"FD", x"20", x"A0", x"E5", x"20", x"44", x"E5", x"A9",
x"00", x"8D", x"19", x"03", x"A2", x"14", x"A0", x"0E",
x"20", x"0C", x"E5", x"A2", x"5C", x"20", x"50", x"F9",
x"68", x"F0", x"17", x"48", x"A2", x"02", x"A0", x"02",
x"20", x"0C", x"E5", x"68", x"48", x"20", x"0D", x"FB",
x"68", x"C9", x"01", x"D0", x"05", x"A2", x"68", x"20",
x"50", x"F9", x"A2", x"00", x"8E", x"20", x"D0", x"E8",
x"10", x"FD", x"A2", x"06", x"8E", x"20", x"D0", x"EA",
x"D0", x"F0", x"A5", x"CC", x"D0", x"43", x"C6", x"CD",
x"10", x"3F", x"A5", x"CF", x"D0", x"27", x"20", x"FC",
x"F8", x"B1", x"D1", x"85", x"CE", x"49", x"80", x"91",
x"D1", x"B1", x"F3", x"8D", x"87", x"02", x"AD", x"86",
x"02", x"91", x"F3", x"A9", x"01", x"85", x"CF", x"D0",
x"1C", x"A9", x"80", x"85", x"CC", x"A9", x"FF", x"85",
x"CD", x"A5", x"CF", x"F0", x"10", x"20", x"FC", x"F8",
x"A5", x"CE", x"91", x"D1", x"AD", x"87", x"02", x"91",
x"F3", x"A9", x"00", x"85", x"CF", x"A9", x"14", x"85",
x"CD", x"60", x"20", x"C5", x"ED", x"A5", x"D7", x"AA",
x"29", x"60", x"D0", x"03", x"4C", x"EE", x"FD", x"8A",
x"20", x"1F", x"E7", x"AA", x"20", x"FC", x"F8", x"8A",
x"05", x"C7", x"91", x"D1", x"A5", x"D8", x"F0", x"02",
x"C6", x"D8", x"8A", x"20", x"09", x"F9", x"AD", x"86",
x"02", x"91", x"F3", x"A4", x"D3", x"C8", x"84", x"D3",
x"C0", x"28", x"D0", x"07", x"20", x"64", x"F6", x"E6",
x"D6", x"A4", x"D3", x"C0", x"50", x"90", x"03", x"4C",
x"BF", x"F9", x"20", x"6C", x"E5", x"20", x"7A", x"F9",
x"4C", x"F1", x"F1", x"A9", x"00", x"85", x"AB", x"85",
x"9F", x"85", x"9E", x"A0", x"89", x"20", x"15", x"EA",
x"B0", x"40", x"20", x"0F", x"FA", x"20", x"74", x"EC",
x"90", x"1C", x"BA", x"E0", x"20", x"90", x"33", x"A6",
x"9E", x"A5", x"C3", x"9D", x"00", x"01", x"E8", x"A5",
x"C4", x"9D", x"00", x"01", x"E8", x"86", x"9E", x"20",
x"0F", x"FA", x"90", x"16", x"B0", x"1A", x"20", x"0F",
x"FA", x"90", x"06", x"20", x"0F", x"F8", x"4C", x"78",
x"EE", x"A5", x"A7", x"A0", x"00", x"91", x"C3", x"20",
x"0F", x"F8", x"20", x"B9", x"FE", x"4C", x"3D", x"EE",
x"18", x"60", x"38", x"60", x"AD", x"00", x"DD", x"09",
x"08", x"8D", x"00", x"DD", x"AD", x"00", x"DD", x"09",
x"10", x"8D", x"00", x"DD", x"29", x"DF", x"D0", x"3A",
x"AD", x"00", x"DD", x"09", x"10", x"D0", x"F5", x"AD",
x"00", x"DD", x"29", x"F7", x"8D", x"00", x"DD", x"AD",
x"00", x"DD", x"29", x"DF", x"8D", x"00", x"DD", x"29",
x"EF", x"4C", x"CA", x"EE", x"AD", x"00", x"DD", x"09",
x"20", x"8D", x"00", x"DD", x"29", x"EF", x"D0", x"12",
x"AD", x"00", x"DD", x"09", x"20", x"8D", x"00", x"DD",
x"29", x"EF", x"8D", x"00", x"DD", x"AD", x"00", x"DD",
x"29", x"F7", x"8D", x"00", x"DD", x"60", x"A0", x"09",
x"20", x"15", x"EA", x"B0", x"34", x"20", x"0F", x"FA",
x"20", x"74", x"EC", x"90", x"02", x"B0", x"1A", x"20",
x"0A", x"EF", x"F0", x"07", x"20", x"0F", x"FA", x"B0",
x"16", x"90", x"0E", x"20", x"0F", x"FA", x"B0", x"06",
x"A5", x"A7", x"A0", x"00", x"91", x"C3", x"20", x"0F",
x"F8", x"20", x"B9", x"FE", x"4C", x"D8", x"EE", x"A5",
x"9E", x"C5", x"9F", x"D0", x"04", x"A5", x"AB", x"C9",
x"01", x"60", x"A6", x"9F", x"BD", x"00", x"01", x"C5",
x"C3", x"D0", x"0D", x"BD", x"01", x"01", x"C5", x"C4",
x"D0", x"06", x"E6", x"9F", x"E6", x"9F", x"A9", x"00",
x"60", x"A5", x"A3", x"C9", x"01", x"D0", x"03", x"4C",
x"6C", x"F1", x"8A", x"48", x"98", x"48", x"78", x"20",
x"6D", x"E9", x"20", x"9F", x"EE", x"20", x"E2", x"F7",
x"20", x"93", x"FA", x"A5", x"A3", x"C9", x"02", x"D0",
x"07", x"AD", x"01", x"DD", x"48", x"4C", x"6E", x"EF",
x"A2", x"07", x"A9", x"00", x"48", x"20", x"6D", x"E9",
x"AD", x"00", x"DD", x"2A", x"10", x"FA", x"68", x"6A",
x"48", x"A0", x"19", x"AD", x"00", x"DD", x"2A", x"10",
x"0A", x"88", x"D0", x"F7", x"20", x"A0", x"F9", x"68",
x"4C", x"74", x"EF", x"CA", x"10", x"DF", x"20", x"AC",
x"EE", x"68", x"85", x"A4", x"68", x"A8", x"68", x"AA",
x"A5", x"A4", x"18", x"58", x"60", x"78", x"AD", x"11",
x"D0", x"85", x"A4", x"20", x"FB", x"F1", x"20", x"17",
x"E7", x"A0", x"FF", x"20", x"6D", x"E9", x"AD", x"00",
x"DD", x"29", x"DF", x"EA", x"20", x"9B", x"F9", x"8D",
x"00", x"DD", x"A5", x"94", x"09", x"20", x"AA", x"EA",
x"EA", x"AD", x"00", x"DD", x"4A", x"4A", x"EA", x"0D",
x"00", x"DD", x"4A", x"4A", x"45", x"94", x"4D", x"00",
x"DD", x"4A", x"4A", x"45", x"94", x"4D", x"00", x"DD",
x"C8", x"91", x"AE", x"2C", x"00", x"DD", x"8E", x"00",
x"DD", x"70", x"09", x"C0", x"FF", x"D0", x"C4", x"E6",
x"AF", x"4C", x"8B", x"EF", x"AA", x"38", x"20", x"76",
x"F8", x"A9", x"00", x"85", x"94", x"A9", x"01", x"85",
x"A3", x"A5", x"A4", x"8D", x"11", x"D0", x"86", x"A4",
x"4C", x"DF", x"E7", x"20", x"4C", x"F0", x"20", x"1A",
x"ED", x"B0", x"08", x"20", x"43", x"F0", x"20", x"2B",
x"EE", x"90", x"06", x"20", x"B0", x"FE", x"4C", x"26",
x"F4", x"20", x"43", x"F0", x"20", x"CE", x"EE", x"B0",
x"F2", x"A0", x"00", x"B1", x"B2", x"C9", x"05", x"D0",
x"03", x"4C", x"B0", x"E6", x"C9", x"01", x"F0", x"08",
x"C9", x"03", x"D0", x"CF", x"A9", x"01", x"85", x"B9",
x"20", x"B0", x"FE", x"20", x"F9", x"E5", x"B0", x"C3",
x"20", x"28", x"ED", x"A0", x"00", x"20", x"2B", x"EE",
x"90", x"03", x"4C", x"B0", x"E6", x"20", x"C0", x"FE",
x"F0", x"03", x"4C", x"B0", x"E6", x"20", x"B0", x"FE",
x"20", x"CE", x"EE", x"90", x"03", x"4C", x"B0", x"E6",
x"4C", x"A7", x"E6", x"A5", x"B3", x"85", x"C4", x"A5",
x"B2", x"85", x"C3", x"60", x"A5", x"C4", x"85", x"C2",
x"A5", x"C3", x"85", x"C1", x"60", x"4C", x"43", x"FF",
x"A5", x"B7", x"D0", x"03", x"4C", x"7F", x"FC", x"20",
x"23", x"FF", x"A5", x"BA", x"20", x"6A", x"F9", x"B0",
x"EC", x"A9", x"01", x"20", x"72", x"E5", x"B0", x"E5",
x"20", x"5C", x"FB", x"B0", x"E0", x"A5", x"BA", x"20",
x"6A", x"F9", x"B0", x"D9", x"A9", x"61", x"85", x"A4",
x"20", x"DA", x"FA", x"B0", x"D0", x"20", x"61", x"FF",
x"A5", x"C1", x"85", x"A4", x"18", x"20", x"C9", x"F0",
x"A5", x"C2", x"85", x"A4", x"18", x"20", x"C9", x"F0",
x"20", x"B0", x"FE", x"A0", x"00", x"20", x"92", x"EB",
x"85", x"A4", x"18", x"20", x"C9", x"F0", x"20", x"B9",
x"FE", x"20", x"C0", x"FE", x"D0", x"EF", x"A5", x"BA",
x"20", x"09", x"FD", x"A5", x"BA", x"20", x"6A", x"F9",
x"A9", x"E1", x"85", x"A4", x"20", x"DA", x"FA", x"20",
x"CD", x"F4", x"A5", x"BA", x"20", x"09", x"FD", x"18",
x"60", x"08", x"A5", x"A3", x"C9", x"01", x"D0", x"04",
x"28", x"4C", x"C8", x"F2", x"28", x"8A", x"48", x"98",
x"48", x"20", x"97", x"EE", x"78", x"20", x"E2", x"F7",
x"90", x"06", x"20", x"E8", x"F7", x"20", x"E2", x"F7",
x"A5", x"A3", x"C9", x"02", x"D0", x"10", x"A9", x"FF",
x"8D", x"03", x"DD", x"A5", x"A4", x"8D", x"01", x"DD",
x"20", x"90", x"EE", x"4C", x"2B", x"F1", x"20", x"90",
x"EE", x"20", x"EE", x"F7", x"A2", x"07", x"D0", x"07",
x"A5", x"A3", x"F0", x"03", x"20", x"F3", x"FA", x"A5",
x"A4", x"4A", x"85", x"A4", x"B0", x"06", x"20", x"AC",
x"EE", x"4C", x"1F", x"F1", x"20", x"9F", x"EE", x"20",
x"FA", x"F7", x"20", x"90", x"EE", x"20", x"FA", x"F7",
x"CA", x"10", x"DB", x"58", x"A2", x"FF", x"AD", x"00",
x"DD", x"10", x"08", x"CA", x"D0", x"F8", x"30", x"03",
x"4C", x"CC", x"FA", x"4C", x"C2", x"FA", x"4C", x"8A",
x"F8", x"2A", x"A5", x"C6", x"D0", x"02", x"38", x"60",
x"AD", x"77", x"02", x"48", x"98", x"48", x"20", x"1D",
x"FD", x"68", x"A8", x"68", x"18", x"60", x"00", x"A5",
x"99", x"D0", x"03", x"4C", x"73", x"E9", x"20", x"1A",
x"F9", x"B0", x"03", x"4C", x"7A", x"FE", x"4C", x"43",
x"FF", x"6C", x"8F", x"02", x"78", x"8A", x"48", x"98",
x"48", x"20", x"CB", x"F8", x"48", x"20", x"6D", x"E9",
x"AD", x"00", x"DD", x"29", x"DF", x"AA", x"20", x"02",
x"E7", x"8E", x"00", x"DD", x"A5", x"94", x"09", x"20",
x"AA", x"EA", x"EA", x"AD", x"00", x"DD", x"4A", x"4A",
x"EA", x"0D", x"00", x"DD", x"4A", x"4A", x"45", x"94",
x"4D", x"00", x"DD", x"4A", x"4A", x"45", x"94", x"4D",
x"00", x"DD", x"85", x"A4", x"EA", x"EA", x"2C", x"00",
x"DD", x"8E", x"00", x"DD", x"50", x"08", x"AD", x"00",
x"DD", x"30", x"12", x"20", x"A0", x"F9", x"A9", x"00",
x"85", x"94", x"A9", x"01", x"85", x"A3", x"68", x"8D",
x"15", x"D0", x"4C", x"74", x"EF", x"20", x"85", x"FC",
x"B0", x"EC", x"85", x"D7", x"8A", x"48", x"98", x"48",
x"08", x"A5", x"9A", x"C9", x"03", x"D0", x"03", x"4C",
x"E2", x"ED", x"20", x"1A", x"F9", x"B0", x"03", x"4C",
x"23", x"F9", x"28", x"68", x"A8", x"68", x"AA", x"38",
x"60", x"28", x"68", x"A8", x"68", x"AA", x"4C", x"43",
x"FF", x"28", x"58", x"68", x"A8", x"68", x"AA", x"A5",
x"D7", x"18", x"60", x"AD", x"11", x"D0", x"29", x"EF",
x"8D", x"11", x"D0", x"AD", x"11", x"D0", x"10", x"FB",
x"AD", x"11", x"D0", x"30", x"FB", x"60", x"48", x"98",
x"48", x"20", x"9C", x"F9", x"8A", x"20", x"3E", x"F9",
x"90", x"03", x"4C", x"90", x"EA", x"B9", x"63", x"02",
x"F0", x"0F", x"20", x"1A", x"F9", x"B0", x"03", x"4C",
x"42", x"FC", x"C9", x"03", x"F0", x"03", x"4C", x"87",
x"EA", x"B9", x"63", x"02", x"85", x"99", x"68", x"A8",
x"68", x"18", x"60", x"68", x"A8", x"68", x"4C", x"79",
x"FC", x"90", x"06", x"AC", x"82", x"02", x"AE", x"81",
x"02", x"8C", x"82", x"02", x"8E", x"81", x"02", x"60",
x"48", x"98", x"48", x"20", x"9C", x"F9", x"8A", x"20",
x"3E", x"F9", x"90", x"03", x"4C", x"90", x"EA", x"B9",
x"63", x"02", x"F0", x"17", x"20", x"1A", x"F9", x"B0",
x"03", x"4C", x"21", x"E5", x"C9", x"03", x"F0", x"03",
x"4C", x"87", x"EA", x"B9", x"63", x"02", x"85", x"9A",
x"4C", x"36", x"F2", x"68", x"A8", x"68", x"4C", x"7C",
x"FC", x"78", x"D8", x"48", x"AD", x"19", x"03", x"F0",
x"04", x"68", x"6C", x"18", x"03", x"68", x"4C", x"47",
x"FE", x"20", x"3E", x"F9", x"B0", x"28", x"B9", x"63",
x"02", x"20", x"1A", x"F9", x"B0", x"03", x"4C", x"FB",
x"F3", x"C8", x"C0", x"0A", x"10", x"15", x"B9", x"59",
x"02", x"99", x"58", x"02", x"B9", x"63", x"02", x"99",
x"62", x"02", x"B9", x"6D", x"02", x"99", x"6C", x"02",
x"4C", x"A1", x"F2", x"C6", x"98", x"18", x"60", x"78",
x"84", x"A0", x"86", x"A1", x"85", x"A2", x"58", x"60",
x"78", x"90", x"02", x"C6", x"A3", x"8A", x"48", x"98",
x"48", x"20", x"C5", x"EE", x"20", x"CB", x"F8", x"48",
x"A5", x"A4", x"29", x"0F", x"AA", x"BD", x"5A", x"F9",
x"48", x"A5", x"A4", x"29", x"F0", x"48", x"A6", x"94",
x"20", x"E2", x"F7", x"20", x"02", x"E7", x"8E", x"00",
x"DD", x"68", x"05", x"94", x"8D", x"00", x"DD", x"4A",
x"4A", x"29", x"30", x"05", x"94", x"8D", x"00", x"DD",
x"68", x"05", x"94", x"8D", x"00", x"DD", x"4A", x"4A",
x"29", x"30", x"8D", x"00", x"DD", x"A5", x"94", x"A6",
x"A3", x"F0", x"11", x"09", x"10", x"8D", x"00", x"DD",
x"A9", x"01", x"85", x"A3", x"68", x"8D", x"15", x"D0",
x"58", x"4C", x"C2", x"FA", x"8D", x"00", x"DD", x"20",
x"FA", x"F7", x"A5", x"94", x"4C", x"13", x"F3", x"4C",
x"AA", x"FA", x"00", x"20", x"E5", x"F9", x"A9", x"00",
x"85", x"99", x"A9", x"03", x"85", x"9A", x"60", x"A2",
x"00", x"86", x"01", x"91", x"C3", x"A2", x"00", x"86",
x"01", x"60", x"20", x"9C", x"F9", x"A4", x"98", x"F0",
x"10", x"88", x"B9", x"59", x"02", x"C5", x"B8", x"D0",
x"03", x"4C", x"6D", x"FC", x"C0", x"00", x"4C", x"4F",
x"F3", x"A4", x"98", x"C0", x"0A", x"90", x"03", x"4C",
x"6A", x"FC", x"A5", x"B8", x"99", x"59", x"02", x"A5",
x"BA", x"99", x"63", x"02", x"A5", x"B9", x"99", x"6D",
x"02", x"C8", x"84", x"98", x"A5", x"BA", x"20", x"1A",
x"F9", x"B0", x"03", x"4C", x"7D", x"FE", x"18", x"60",
x"09", x"90", x"4C", x"DA", x"F9", x"A6", x"D8", x"F0",
x"05", x"A9", x"14", x"4C", x"80", x"F8", x"A4", x"D3",
x"F0", x"47", x"C0", x"28", x"D0", x"16", x"A5", x"F3",
x"D0", x"04", x"C6", x"F4", x"C6", x"D2", x"C6", x"F3",
x"C6", x"D1", x"A2", x"27", x"A0", x"00", x"20", x"CC",
x"F3", x"4C", x"CE", x"EC", x"20", x"FC", x"F8", x"84",
x"D3", x"20", x"50", x"FA", x"98", x"38", x"E5", x"D3",
x"AA", x"A4", x"D3", x"88", x"20", x"CC", x"F3", x"C6",
x"D3", x"4C", x"22", x"EE", x"C8", x"B1", x"F3", x"88",
x"91", x"F3", x"C8", x"B1", x"D1", x"88", x"91", x"D1",
x"C8", x"CA", x"10", x"F0", x"A9", x"20", x"91", x"D1",
x"60", x"A4", x"D6", x"F0", x"E4", x"C6", x"D6", x"A9",
x"27", x"85", x"D3", x"20", x"E6", x"EB", x"A0", x"27",
x"A9", x"20", x"91", x"D1", x"D0", x"D3", x"60", x"3C",
x"02", x"07", x"00", x"20", x"B5", x"F8", x"B9", x"6D",
x"02", x"C9", x"60", x"D0", x"06", x"20", x"24", x"FA",
x"4C", x"A1", x"F2", x"05", x"E0", x"85", x"A4", x"20",
x"DA", x"FA", x"B0", x"03", x"20", x"CD", x"F4", x"4C",
x"A1", x"F2", x"20", x"62", x"F8", x"20", x"C0", x"F8",
x"20", x"7C", x"FA", x"20", x"D4", x"E5", x"20", x"96",
x"EA", x"B0", x"03", x"4C", x"E3", x"EF", x"20", x"E0",
x"EC", x"90", x"03", x"4C", x"E3", x"EF", x"A0", x"00",
x"91", x"B2", x"C8", x"20", x"5A", x"E9", x"91", x"B2",
x"C8", x"C0", x"05", x"D0", x"03", x"20", x"5A", x"E9",
x"C0", x"C0", x"D0", x"EF", x"A0", x"00", x"B1", x"B2",
x"F0", x"08", x"29", x"01", x"D0", x"04", x"A9", x"01",
x"85", x"B9", x"20", x"C0", x"F8", x"20", x"F9", x"E5",
x"B0", x"CC", x"A2", x"0A", x"BD", x"3F", x"F3", x"9D",
x"00", x"01", x"CA", x"10", x"F7", x"A5", x"01", x"8D",
x"07", x"01", x"A9", x"00", x"85", x"9B", x"20", x"FE",
x"EC", x"B0", x"FB", x"20", x"5A", x"E9", x"20", x"00",
x"01", x"45", x"9B", x"85", x"9B", x"20", x"B9", x"FE",
x"20", x"C0", x"FE", x"D0", x"EE", x"20", x"5A", x"E9",
x"AA", x"20", x"C0", x"F8", x"E4", x"9B", x"D0", x"03",
x"4C", x"A7", x"E6", x"4C", x"B0", x"E6", x"84", x"C4",
x"86", x"C3", x"6C", x"30", x"03", x"85", x"93", x"A5",
x"C3", x"85", x"C1", x"A5", x"C4", x"84", x"C2", x"20",
x"9C", x"F9", x"A5", x"BA", x"C9", x"01", x"D0", x"03",
x"4C", x"1A", x"F4", x"C9", x"07", x"D0", x"03", x"4C",
x"1A", x"F4", x"20", x"16", x"F9", x"B0", x"03", x"4C",
x"54", x"E7", x"4C", x"49", x"FF", x"8A", x"48", x"98",
x"48", x"20", x"FA", x"F7", x"20", x"AA", x"F8", x"20",
x"FA", x"F7", x"4C", x"C2", x"FA", x"14", x"0D", x"1D",
x"88", x"85", x"86", x"87", x"11", x"33", x"57", x"41",
x"34", x"5A", x"53", x"45", x"00", x"35", x"52", x"44",
x"36", x"43", x"46", x"54", x"58", x"37", x"59", x"47",
x"38", x"42", x"48", x"55", x"56", x"39", x"49", x"4A",
x"30", x"4D", x"4B", x"4F", x"4E", x"2B", x"50", x"4C",
x"2D", x"2E", x"3A", x"40", x"2C", x"5C", x"2A", x"3B",
x"13", x"00", x"3D", x"5E", x"2F", x"31", x"5F", x"00",
x"32", x"20", x"00", x"51", x"03", x"94", x"8D", x"9D",
x"8C", x"89", x"8A", x"8B", x"91", x"23", x"77", x"61",
x"24", x"7A", x"73", x"65", x"00", x"25", x"72", x"64",
x"26", x"63", x"66", x"74", x"78", x"27", x"79", x"67",
x"28", x"62", x"68", x"75", x"76", x"29", x"69", x"6A",
x"92", x"6D", x"6B", x"6F", x"6E", x"DB", x"70", x"6C",
x"DD", x"3E", x"5B", x"BA", x"3C", x"A9", x"C0", x"5D",
x"93", x"00", x"3D", x"DE", x"3F", x"21", x"5F", x"00",
x"22", x"A0", x"00", x"71", x"83", x"94", x"8D", x"9D",
x"8C", x"89", x"8A", x"8B", x"91", x"96", x"B3", x"B0",
x"97", x"AD", x"AE", x"B1", x"00", x"98", x"B2", x"AC",
x"99", x"BC", x"BB", x"A3", x"BD", x"9A", x"B7", x"A5",
x"9B", x"BF", x"B4", x"B8", x"BE", x"30", x"A2", x"B5",
x"30", x"A7", x"A1", x"B9", x"AA", x"A6", x"AF", x"B6",
x"DC", x"3E", x"5B", x"A4", x"3C", x"A8", x"DF", x"5D",
x"93", x"00", x"3D", x"DE", x"3F", x"81", x"5F", x"00",
x"95", x"A0", x"00", x"AB", x"83", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"1C", x"17", x"01",
x"9F", x"1A", x"13", x"05", x"00", x"9C", x"12", x"04",
x"1E", x"03", x"06", x"14", x"18", x"1F", x"19", x"07",
x"9E", x"02", x"08", x"15", x"16", x"12", x"09", x"0A",
x"92", x"0D", x"0B", x"0F", x"0E", x"00", x"10", x"0C",
x"00", x"00", x"1B", x"00", x"00", x"1C", x"00", x"1D",
x"00", x"00", x"1F", x"1E", x"00", x"90", x"06", x"00",
x"05", x"00", x"00", x"11", x"00", x"84", x"AF", x"86",
x"AE", x"AA", x"B5", x"01", x"85", x"C2", x"B5", x"00",
x"85", x"C1", x"6C", x"32", x"03", x"20", x"9C", x"F9",
x"A5", x"BA", x"20", x"16", x"F9", x"B0", x"03", x"4C",
x"58", x"F0", x"4C", x"49", x"FF", x"20", x"1E", x"F8",
x"F0", x"05", x"F0", x"03", x"4C", x"25", x"EE", x"20",
x"50", x"FA", x"A6", x"D6", x"B5", x"D9", x"10", x"12",
x"20", x"32", x"F6", x"A9", x"20", x"91", x"D1", x"20",
x"1E", x"F8", x"F0", x"03", x"20", x"64", x"F6", x"4C",
x"22", x"EE", x"A5", x"D3", x"38", x"E9", x"28", x"85",
x"D3", x"20", x"32", x"F6", x"A9", x"20", x"91", x"D1",
x"D0", x"ED", x"88", x"B1", x"F3", x"C8", x"91", x"F3",
x"88", x"B1", x"D1", x"C8", x"91", x"D1", x"88", x"C4",
x"D3", x"D0", x"EF", x"E6", x"D8", x"60", x"60", x"48",
x"A5", x"94", x"D0", x"07", x"E6", x"94", x"18", x"68",
x"85", x"95", x"60", x"18", x"20", x"C9", x"F0", x"E6",
x"94", x"4C", x"4F", x"F6", x"E6", x"D6", x"4C", x"E6",
x"EB", x"20", x"EA", x"E8", x"A4", x"D6", x"B9", x"D9",
x"00", x"10", x"F1", x"C0", x"18", x"F0", x"F2", x"B9",
x"DA", x"00", x"10", x"EA", x"20", x"FA", x"F9", x"A0",
x"17", x"C4", x"D6", x"F0", x"0B", x"90", x"09", x"B9",
x"D9", x"00", x"99", x"DA", x"00", x"88", x"D0", x"F1",
x"A4", x"D6", x"A9", x"00", x"99", x"DA", x"00", x"A9",
x"17", x"38", x"E5", x"D6", x"F0", x"4B", x"AA", x"AD",
x"88", x"02", x"18", x"69", x"03", x"85", x"AD", x"85",
x"AF", x"A9", x"DB", x"85", x"D2", x"85", x"F4", x"A9",
x"C0", x"85", x"AE", x"85", x"F3", x"A9", x"98", x"85",
x"AC", x"85", x"D1", x"A0", x"27", x"B1", x"AC", x"91",
x"AE", x"B1", x"D1", x"91", x"F3", x"88", x"10", x"F5",
x"A5", x"AC", x"38", x"E9", x"28", x"85", x"AC", x"85",
x"D1", x"B0", x"04", x"C6", x"AD", x"C6", x"D2", x"A5",
x"AE", x"38", x"E9", x"28", x"85", x"AE", x"85", x"F3",
x"B0", x"04", x"C6", x"AF", x"C6", x"F4", x"CA", x"D0",
x"D2", x"20", x"34", x"FE", x"A6", x"D6", x"E8", x"20",
x"FF", x"E9", x"4C", x"B6", x"FC", x"A5", x"91", x"10",
x"04", x"A9", x"FF", x"18", x"60", x"38", x"A9", x"00",
x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"C3", x"C2", x"CD", x"38", x"30", x"A9", x"00", x"85",
x"CC", x"60", x"A9", x"0D", x"4C", x"D2", x"FF", x"A9",
x"20", x"4C", x"D2", x"FF", x"A2", x"FF", x"8E", x"00",
x"DC", x"60", x"AD", x"00", x"DD", x"10", x"FB", x"60",
x"AD", x"00", x"DD", x"30", x"FB", x"60", x"A2", x"0A",
x"CA", x"10", x"FD", x"60", x"20", x"66", x"E5", x"4C",
x"22", x"EE", x"0D", x"FF", x"03", x"0D", x"FF", x"03",
x"60", x"85", x"B8", x"84", x"B9", x"86", x"BA", x"60",
x"85", x"B7", x"84", x"BC", x"86", x"BB", x"60", x"A5",
x"A7", x"45", x"AB", x"85", x"AB", x"60", x"FE", x"FD",
x"FB", x"F7", x"EF", x"DF", x"BF", x"7F", x"20", x"50",
x"FA", x"B1", x"D1", x"C9", x"20", x"60", x"00", x"08",
x"10", x"18", x"20", x"28", x"30", x"38", x"00", x"40",
x"80", x"FF", x"C0", x"FF", x"FF", x"FF", x"00", x"80",
x"00", x"00", x"00", x"00", x"10", x"24", x"A9", x"00",
x"85", x"D4", x"85", x"D8", x"4C", x"25", x"EE", x"78",
x"A4", x"A0", x"A6", x"A1", x"A5", x"A2", x"58", x"60",
x"AD", x"11", x"D0", x"09", x"10", x"8D", x"11", x"D0",
x"60", x"A6", x"BA", x"E0", x"08", x"B0", x"02", x"A2",
x"08", x"60", x"A5", x"93", x"D0", x"01", x"60", x"68",
x"68", x"4C", x"43", x"FF", x"A9", x"80", x"2C", x"A9",
x"00", x"85", x"C7", x"4C", x"25", x"EE", x"98", x"65",
x"AE", x"85", x"AE", x"90", x"02", x"E6", x"AF", x"60",
x"18", x"69", x"80", x"90", x"02", x"69", x"BF", x"4C",
x"F3", x"ED", x"A5", x"99", x"D0", x"03", x"4C", x"42",
x"F1", x"4C", x"5E", x"F1", x"A5", x"90", x"F0", x"04",
x"18", x"A9", x"0D", x"60", x"4C", x"21", x"EF", x"A9",
x"00", x"2C", x"A9", x"80", x"8D", x"91", x"02", x"4C",
x"25", x"EE", x"AD", x"00", x"DD", x"09", x"10", x"29",
x"D7", x"8D", x"00", x"DD", x"60", x"48", x"A5", x"94",
x"F0", x"04", x"38", x"20", x"D5", x"F0", x"68", x"60",
x"A9", x"00", x"A0", x"1C", x"99", x"00", x"D4", x"88",
x"10", x"FA", x"60", x"20", x"17", x"E7", x"AD", x"15",
x"D0", x"A2", x"00", x"8E", x"15", x"D0", x"60", x"FD",
x"BF", x"7F", x"7F", x"80", x"10", x"20", x"04", x"01",
x"01", x"02", x"04", x"A5", x"BA", x"C9", x"02", x"D0",
x"03", x"A9", x"FF", x"60", x"A5", x"90", x"60", x"A5",
x"01", x"09", x"20", x"D0", x"04", x"A5", x"01", x"29",
x"DF", x"85", x"01", x"60", x"A4", x"D3", x"C0", x"28",
x"90", x"04", x"98", x"E9", x"28", x"A8", x"C0", x"00",
x"60", x"C9", x"22", x"D0", x"08", x"A5", x"D4", x"49",
x"80", x"85", x"D4", x"A9", x"22", x"60", x"C9", x"08",
x"90", x"07", x"C9", x"04", x"90", x"03", x"C9", x"1F",
x"60", x"38", x"60", x"A5", x"D7", x"20", x"A8", x"FF",
x"B0", x"03", x"4C", x"F1", x"F1", x"4C", x"E2", x"F1",
x"A2", x"05", x"BD", x"03", x"80", x"DD", x"C7", x"F7",
x"D0", x"03", x"CA", x"D0", x"F5", x"60", x"A4", x"98",
x"88", x"30", x"07", x"D9", x"59", x"02", x"D0", x"F8",
x"18", x"60", x"38", x"60", x"20", x"D2", x"FF", x"E8",
x"BD", x"D1", x"EA", x"10", x"F7", x"29", x"7F", x"4C",
x"D2", x"FF", x"00", x"80", x"20", x"A0", x"40", x"C0",
x"60", x"E0", x"10", x"90", x"30", x"B0", x"50", x"D0",
x"70", x"F0", x"20", x"B5", x"F8", x"20", x"1A", x"F9",
x"90", x"03", x"4C", x"76", x"FC", x"09", x"20", x"4C",
x"73", x"FA", x"A5", x"CC", x"D0", x"0C", x"A5", x"CF",
x"D0", x"08", x"A9", x"01", x"85", x"CD", x"A9", x"00",
x"85", x"CF", x"60", x"A2", x"12", x"AD", x"12", x"D0",
x"CD", x"12", x"D0", x"F0", x"FB", x"AD", x"12", x"D0",
x"CA", x"D0", x"F5", x"60", x"A9", x"00", x"F0", x"0A",
x"A5", x"90", x"09", x"40", x"D0", x"04", x"A5", x"90",
x"09", x"80", x"85", x"90", x"60", x"AD", x"18", x"D0",
x"29", x"02", x"8D", x"18", x"D0", x"4C", x"25", x"EE",
x"AD", x"18", x"D0", x"09", x"02", x"D0", x"F3", x"A4",
x"D6", x"C0", x"18", x"D0", x"03", x"20", x"EA", x"E8",
x"E6", x"D6", x"A9", x"00", x"85", x"D3", x"4C", x"22",
x"EE", x"20", x"B5", x"F8", x"A9", x"FF", x"85", x"A3",
x"A9", x"5F", x"85", x"A4", x"20", x"DA", x"FA", x"B0",
x"03", x"4C", x"AD", x"FB", x"60", x"A5", x"99", x"20",
x"1A", x"F9", x"B0", x"03", x"20", x"D1", x"F9", x"A5",
x"9A", x"20", x"1A", x"F9", x"B0", x"03", x"4C", x"09",
x"FD", x"60", x"68", x"AA", x"68", x"A8", x"A5", x"AC",
x"48", x"A5", x"AE", x"48", x"A5", x"AD", x"48", x"A5",
x"AF", x"48", x"98", x"48", x"8A", x"48", x"60", x"20",
x"91", x"FD", x"C5", x"96", x"B0", x"F9", x"4C", x"91",
x"FD", x"20", x"91", x"FD", x"B0", x"FB", x"C5", x"96",
x"B0", x"F7", x"90", x"F2", x"AA", x"20", x"D1", x"F9",
x"8A", x"20", x"6A", x"F9", x"A9", x"E0", x"85", x"A4",
x"20", x"DA", x"FA", x"20", x"CD", x"F4", x"20", x"09",
x"FD", x"60", x"8A", x"48", x"98", x"48", x"08", x"78",
x"20", x"C5", x"EE", x"20", x"9F", x"EE", x"20", x"6D",
x"E9", x"20", x"84", x"EE", x"28", x"4C", x"C2", x"FA",
x"A4", x"D6", x"C0", x"18", x"B0", x"0D", x"B9", x"D9",
x"00", x"10", x"08", x"B9", x"DA", x"00", x"30", x"03",
x"A0", x"4F", x"60", x"A0", x"27", x"60", x"20", x"B5",
x"F8", x"20", x"1A", x"F9", x"90", x"03", x"4C", x"76",
x"FC", x"09", x"40", x"85", x"A4", x"A9", x"FF", x"85",
x"A3", x"4C", x"DA", x"FA", x"A2", x"03", x"8E", x"04",
x"DD", x"A2", x"00", x"8E", x"05", x"DD", x"8E", x"07",
x"DD", x"CA", x"8E", x"06", x"DD", x"A2", x"11", x"8E",
x"0E", x"DD", x"60", x"A2", x"13", x"2C", x"00", x"DD",
x"50", x"0F", x"CA", x"D0", x"F8", x"20", x"A0", x"F9",
x"20", x"AC", x"EE", x"20", x"EE", x"F7", x"20", x"9F",
x"EE", x"60", x"98", x"48", x"A4", x"98", x"F0", x"0A",
x"88", x"B9", x"59", x"02", x"20", x"C3", x"FF", x"4C",
x"AC", x"FA", x"68", x"A8", x"20", x"33", x"F3", x"4C",
x"9C", x"F9", x"A9", x"00", x"85", x"94", x"68", x"A8",
x"68", x"AA", x"18", x"60", x"20", x"AA", x"F8", x"A9",
x"00", x"85", x"94", x"68", x"A8", x"68", x"AA", x"4C",
x"76", x"FC", x"8A", x"48", x"98", x"48", x"20", x"7C",
x"EE", x"20", x"8B", x"F9", x"AD", x"00", x"DD", x"10",
x"03", x"4C", x"CC", x"FA", x"20", x"9F", x"EE", x"18",
x"4C", x"DC", x"F0", x"A0", x"25", x"AD", x"00", x"DD",
x"10", x"0B", x"88", x"D0", x"F8", x"A5", x"A3", x"10",
x"0B", x"A9", x"00", x"F0", x"05", x"20", x"E2", x"F7",
x"A9", x"01", x"85", x"A3", x"60", x"F8", x"48", x"4A",
x"4A", x"4A", x"4A", x"C9", x"0A", x"69", x"30", x"D8",
x"20", x"D2", x"FF", x"F8", x"68", x"29", x"0F", x"C9",
x"0A", x"69", x"30", x"D8", x"4C", x"D2", x"FF", x"A0",
x"00", x"20", x"41", x"FB", x"26", x"A7", x"A5", x"A7",
x"C9", x"FF", x"D0", x"05", x"C8", x"10", x"F2", x"30",
x"06", x"C9", x"02", x"D0", x"EA", x"18", x"60", x"38",
x"60", x"20", x"91", x"FD", x"B0", x"0C", x"A9", x"01",
x"8D", x"18", x"D4", x"A9", x"06", x"8D", x"20", x"D0",
x"38", x"60", x"A9", x"00", x"8D", x"18", x"D4", x"8D",
x"20", x"D0", x"18", x"60", x"A0", x"00", x"C4", x"B7",
x"F0", x"12", x"20", x"A1", x"EB", x"C8", x"C4", x"B7",
x"18", x"D0", x"01", x"38", x"85", x"A4", x"20", x"C9",
x"F0", x"4C", x"5E", x"FB", x"4C", x"09", x"FD", x"A9",
x"00", x"85", x"D4", x"85", x"D8", x"85", x"C7", x"A4",
x"D6", x"C0", x"18", x"F0", x"0A", x"B9", x"DA", x"00",
x"30", x"05", x"E6", x"D6", x"20", x"E6", x"EB", x"4C",
x"BF", x"F9", x"20", x"EF", x"F8", x"A5", x"9C", x"8D",
x"20", x"D0", x"4C", x"50", x"F8", x"78", x"A9", x"00",
x"85", x"C6", x"AD", x"20", x"D0", x"85", x"9C", x"20",
x"FB", x"F1", x"4C", x"F5", x"F8", x"8A", x"48", x"98",
x"48", x"08", x"78", x"20", x"B8", x"EE", x"A2", x"FF",
x"AD", x"00", x"DD", x"2A", x"10", x"07", x"CA", x"D0",
x"F7", x"28", x"4C", x"CC", x"FA", x"28", x"4C", x"C2",
x"FA", x"A2", x"06", x"DD", x"B9", x"EB", x"F0", x"05",
x"CA", x"10", x"F8", x"38", x"60", x"BD", x"DF", x"EB",
x"AA", x"BD", x"C0", x"EB", x"F0", x"06", x"20", x"CA",
x"F1", x"E8", x"D0", x"F5", x"18", x"60", x"20", x"91",
x"FD", x"90", x"0C", x"20", x"91", x"FD", x"B0", x"11",
x"A9", x"00", x"8D", x"20", x"D0", x"18", x"60", x"20",
x"91", x"FD", x"90", x"05", x"18", x"A9", x"06", x"D0",
x"F1", x"38", x"60", x"84", x"C4", x"86", x"C3", x"A9",
x"00", x"8D", x"19", x"03", x"A0", x"1F", x"90", x"07",
x"B9", x"14", x"03", x"91", x"C3", x"B0", x"05", x"B1",
x"C3", x"99", x"14", x"03", x"88", x"10", x"F8", x"60",
x"A9", x"48", x"8D", x"8F", x"02", x"A9", x"EB", x"8D",
x"90", x"02", x"A9", x"01", x"85", x"CD", x"85", x"CC",
x"A2", x"01", x"8E", x"86", x"02", x"A2", x"0A", x"8E",
x"89", x"02", x"A2", x"00", x"8E", x"91", x"02", x"4C",
x"44", x"E5", x"B9", x"59", x"02", x"C9", x"01", x"D0",
x"03", x"4C", x"3B", x"F2", x"B9", x"63", x"02", x"20",
x"66", x"FA", x"90", x"03", x"4C", x"87", x"EA", x"B9",
x"59", x"02", x"09", x"60", x"20", x"88", x"F3", x"90",
x"03", x"4C", x"87", x"EA", x"4C", x"31", x"F2", x"A9",
x"00", x"2C", x"A9", x"01", x"2C", x"A9", x"02", x"2C",
x"A9", x"03", x"2C", x"A9", x"04", x"2C", x"A9", x"05",
x"2C", x"A9", x"06", x"2C", x"A9", x"07", x"2C", x"A9",
x"08", x"2C", x"A9", x"09", x"2C", x"A9", x"02", x"2C",
x"A9", x"F0", x"38", x"60", x"AD", x"12", x"D0", x"CD",
x"12", x"D0", x"F0", x"FB", x"30", x"F6", x"C9", x"07",
x"90", x"03", x"A9", x"01", x"2C", x"A9", x"00", x"8D",
x"A6", x"02", x"AE", x"A6", x"02", x"F0", x"02", x"A2",
x"01", x"BD", x"F8", x"FF", x"8D", x"04", x"DC", x"BD",
x"EC", x"FD", x"8D", x"05", x"DC", x"60", x"A4", x"D6",
x"B9", x"D9", x"00", x"08", x"20", x"FC", x"F8", x"28",
x"30", x"05", x"98", x"18", x"69", x"28", x"A8", x"84",
x"D3", x"A4", x"D6", x"B9", x"D9", x"00", x"10", x"0D",
x"C0", x"18", x"F0", x"06", x"C8", x"B9", x"D9", x"00",
x"10", x"03", x"A9", x"27", x"2C", x"A9", x"4F", x"85",
x"D5", x"60", x"78", x"D8", x"A9", x"00", x"8D", x"19",
x"03", x"A2", x"FF", x"9A", x"20", x"30", x"F9", x"D0",
x"03", x"6C", x"00", x"80", x"A2", x"28", x"8E", x"16",
x"D0", x"20", x"84", x"FF", x"20", x"87", x"FF", x"20",
x"8A", x"FF", x"20", x"81", x"FF", x"58", x"6C", x"00",
x"A0", x"20", x"B5", x"F8", x"A9", x"FF", x"85", x"A3",
x"A9", x"3F", x"4C", x"89", x"E5", x"18", x"A0", x"FD",
x"A2", x"30", x"4C", x"03", x"FC", x"A0", x"01", x"78",
x"B9", x"77", x"02", x"99", x"76", x"02", x"C8", x"CC",
x"89", x"02", x"D0", x"F4", x"C6", x"C6", x"58", x"60",
x"31", x"EA", x"66", x"FE", x"47", x"FE", x"4A", x"F3",
x"91", x"F2", x"0E", x"F2", x"50", x"F2", x"33", x"F3",
x"57", x"F1", x"CA", x"F1", x"ED", x"F6", x"3E", x"F1",
x"2F", x"F3", x"66", x"FE", x"A5", x"F4", x"ED", x"F5",
x"A0", x"00", x"A9", x"00", x"99", x"00", x"03", x"99",
x"00", x"02", x"99", x"02", x"00", x"C8", x"D0", x"F4",
x"A2", x"3C", x"86", x"B2", x"A2", x"03", x"86", x"B3",
x"A2", x"04", x"8E", x"88", x"02", x"A2", x"08", x"8E",
x"82", x"02", x"AE", x"00", x"80", x"E8", x"8E", x"00",
x"80", x"EC", x"00", x"80", x"D0", x"0A", x"A0", x"A0",
x"8C", x"84", x"02", x"CA", x"8E", x"00", x"80", x"60",
x"A0", x"80", x"D0", x"F4", x"8D", x"85", x"02", x"60",
x"60", x"A9", x"10", x"2C", x"0D", x"DC", x"F0", x"FB",
x"AD", x"06", x"DD", x"A2", x"51", x"8E", x"0F", x"DD",
x"C5", x"92", x"60", x"A2", x"27", x"86", x"01", x"A2",
x"2F", x"86", x"00", x"A2", x"7F", x"8E", x"0D", x"DC",
x"8E", x"0D", x"DD", x"8E", x"00", x"DC", x"A9", x"00",
x"8D", x"18", x"D4", x"A2", x"FF", x"8E", x"02", x"DC",
x"E8", x"8E", x"03", x"DC", x"8E", x"03", x"DD", x"A9",
x"3F", x"8D", x"02", x"DD", x"A2", x"08", x"8E", x"0F",
x"DC", x"8E", x"0E", x"DD", x"8E", x"0F", x"DD", x"A2",
x"07", x"8E", x"00", x"DD", x"20", x"A2", x"FC", x"A2",
x"11", x"8E", x"0E", x"DC", x"A2", x"81", x"8E", x"0D",
x"DC", x"4C", x"AA", x"F8", x"42", x"40", x"8A", x"A2",
x"0F", x"E0", x"0C", x"D0", x"0C", x"A8", x"A5", x"D4",
x"05", x"D8", x"F0", x"04", x"98", x"4C", x"80", x"F8",
x"98", x"DD", x"13", x"EC", x"D0", x"09", x"BD", x"33",
x"EC", x"48", x"BD", x"23", x"EC", x"48", x"60", x"CA",
x"10", x"DF", x"A2", x"0F", x"DD", x"DA", x"E8", x"D0",
x"06", x"8E", x"86", x"02", x"4C", x"25", x"EE", x"CA",
x"10", x"F2", x"4C", x"25", x"EE", x"90", x"06", x"AC",
x"84", x"02", x"AE", x"83", x"02", x"8C", x"84", x"02",
x"8E", x"83", x"02", x"60", x"68", x"AA", x"68", x"A8",
x"68", x"85", x"AF", x"68", x"85", x"AD", x"68", x"85",
x"AE", x"68", x"85", x"AC", x"4C", x"0A", x"FA", x"48",
x"8A", x"48", x"98", x"48", x"20", x"30", x"F9", x"D0",
x"03", x"6C", x"02", x"80", x"20", x"E1", x"FF", x"B0",
x"03", x"4C", x"81", x"EA", x"A9", x"00", x"85", x"B0",
x"85", x"B1", x"6C", x"16", x"03", x"00", x"78", x"A2",
x"00", x"8D", x"16", x"D0", x"D8", x"20", x"8A", x"FF",
x"20", x"84", x"FF", x"20", x"5B", x"FF", x"58", x"6C",
x"02", x"A0", x"4C", x"A5", x"FF", x"A4", x"B7", x"F0",
x"15", x"20", x"6A", x"F9", x"90", x"03", x"4C", x"76",
x"FC", x"A5", x"B9", x"20", x"72", x"E5", x"90", x"03",
x"4C", x"76", x"FC", x"20", x"5C", x"FB", x"4C", x"86",
x"F3", x"A4", x"93", x"D0", x"06", x"A0", x"00", x"91",
x"AE", x"18", x"60", x"85", x"A4", x"A0", x"00", x"20",
x"AD", x"EB", x"C5", x"A4", x"F0", x"F3", x"38", x"60",
x"A5", x"C1", x"85", x"C3", x"A5", x"C2", x"85", x"C4",
x"60", x"E6", x"C3", x"D0", x"02", x"E6", x"C4", x"60",
x"A5", x"C4", x"C5", x"AF", x"D0", x"04", x"A5", x"C3",
x"C5", x"AE", x"60", x"A5", x"9D", x"10", x"15", x"A2",
x"00", x"20", x"50", x"F9", x"A0", x"00", x"C4", x"B7",
x"F0", x"0A", x"20", x"A1", x"EB", x"20", x"D2", x"FF",
x"C8", x"4C", x"D6", x"FE", x"60", x"A5", x"9D", x"10",
x"FB", x"A2", x"0F", x"A5", x"93", x"F0", x"02", x"A2",
x"17", x"20", x"50", x"F9", x"A2", x"29", x"20", x"50",
x"F9", x"A5", x"BA", x"C9", x"01", x"F0", x"0E", x"C9",
x"07", x"F0", x"0A", x"A5", x"AF", x"20", x"0D", x"FB",
x"A5", x"AE", x"4C", x"0D", x"FB", x"A5", x"C2", x"20",
x"0D", x"FB", x"A5", x"C1", x"4C", x"0D", x"FB", x"A5",
x"9D", x"10", x"C9", x"A2", x"30", x"20", x"50", x"F9",
x"4C", x"03", x"FF", x"A5", x"9D", x"10", x"BD", x"A2",
x"21", x"20", x"50", x"F9", x"A0", x"00", x"C4", x"B7",
x"F0", x"08", x"B1", x"BB", x"20", x"D2", x"FF", x"C8",
x"D0", x"F4", x"60", x"38", x"60", x"A6", x"AE", x"A4",
x"AF", x"18", x"60", x"20", x"A6", x"F9", x"4C", x"76",
x"FC", x"20", x"A6", x"F9", x"4C", x"82", x"FC", x"A5",
x"93", x"D0", x"04", x"A9", x"1D", x"D0", x"E4", x"A9",
x"1C", x"38", x"60", x"20", x"18", x"E5", x"4C", x"8C",
x"FC", x"A9", x"7F", x"8D", x"0D", x"DD", x"A9", x"00",
x"8D", x"03", x"DD", x"A2", x"20", x"AD", x"0D", x"DD",
x"C9", x"10", x"F0", x"07", x"AD", x"01", x"DD", x"CA",
x"D0", x"F3", x"60", x"A9", x"02", x"85", x"A3", x"60",
x"F0", x"4C", x"5B", x"FF", x"4C", x"A3", x"FD", x"4C",
x"50", x"FD", x"4C", x"15", x"FD", x"4C", x"1A", x"FD",
x"4C", x"1E", x"E5", x"4C", x"B7", x"E6", x"4C", x"88",
x"F3", x"4C", x"25", x"FE", x"4C", x"41", x"F2", x"4C",
x"FD", x"E7", x"4C", x"8C", x"FD", x"4C", x"94", x"F8",
x"4C", x"47", x"F6", x"4C", x"D1", x"F9", x"4C", x"09",
x"FD", x"4C", x"6A", x"F9", x"4C", x"66", x"FA", x"4C",
x"E3", x"F8", x"4C", x"01", x"F8", x"4C", x"08", x"F8",
x"6C", x"1A", x"03", x"6C", x"1C", x"03", x"6C", x"1E",
x"03", x"6C", x"20", x"03", x"6C", x"22", x"03", x"6C",
x"24", x"03", x"6C", x"26", x"03", x"4C", x"9E", x"F4",
x"4C", x"DD", x"F5", x"4C", x"BF", x"F2", x"4C", x"47",
x"F8", x"6C", x"28", x"03", x"6C", x"2A", x"03", x"6C",
x"2C", x"03", x"4C", x"D3", x"E4", x"4C", x"C9", x"E5",
x"4C", x"0A", x"E5", x"A0", x"DC", x"A2", x"00", x"60",
x"95", x"25", x"81", x"F2", x"E2", x"FC", x"53", x"EA"
);
end rom_kernal_pack;
